VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO W_IO
  CLASS BLOCK ;
  FOREIGN W_IO ;
  ORIGIN 0.000 0.000 ;
  SIZE 110.000 BY 390.000 ;
  PIN A_I_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1.400 2.000 1.960 ;
    END
  END A_I_top
  PIN A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 18.200 2.000 18.760 ;
    END
  END A_O_top
  PIN A_T_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 9.240 2.000 9.800 ;
    END
  END A_T_top
  PIN A_config_C_bit0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 51.800 2.000 52.360 ;
    END
  END A_config_C_bit0
  PIN A_config_C_bit1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 59.640 2.000 60.200 ;
    END
  END A_config_C_bit1
  PIN A_config_C_bit2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 68.600 2.000 69.160 ;
    END
  END A_config_C_bit2
  PIN A_config_C_bit3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 76.440 2.000 77.000 ;
    END
  END A_config_C_bit3
  PIN B_I_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 26.040 2.000 26.600 ;
    END
  END B_I_top
  PIN B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 42.840 2.000 43.400 ;
    END
  END B_O_top
  PIN B_T_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 35.000 2.000 35.560 ;
    END
  END B_T_top
  PIN B_config_C_bit0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 85.400 2.000 85.960 ;
    END
  END B_config_C_bit0
  PIN B_config_C_bit1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 93.240 2.000 93.800 ;
    END
  END B_config_C_bit1
  PIN B_config_C_bit2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 102.200 2.000 102.760 ;
    END
  END B_config_C_bit2
  PIN B_config_C_bit3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 111.160 2.000 111.720 ;
    END
  END B_config_C_bit3
  PIN E1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 1.400 110.000 1.960 ;
    END
  END E1BEG[0]
  PIN E1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 3.640 110.000 4.200 ;
    END
  END E1BEG[1]
  PIN E1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 7.000 110.000 7.560 ;
    END
  END E1BEG[2]
  PIN E1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 10.360 110.000 10.920 ;
    END
  END E1BEG[3]
  PIN E2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 12.600 110.000 13.160 ;
    END
  END E2BEG[0]
  PIN E2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 15.960 110.000 16.520 ;
    END
  END E2BEG[1]
  PIN E2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 19.320 110.000 19.880 ;
    END
  END E2BEG[2]
  PIN E2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 21.560 110.000 22.120 ;
    END
  END E2BEG[3]
  PIN E2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 24.920 110.000 25.480 ;
    END
  END E2BEG[4]
  PIN E2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 28.280 110.000 28.840 ;
    END
  END E2BEG[5]
  PIN E2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 31.640 110.000 32.200 ;
    END
  END E2BEG[6]
  PIN E2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 33.880 110.000 34.440 ;
    END
  END E2BEG[7]
  PIN E2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 37.240 110.000 37.800 ;
    END
  END E2BEGb[0]
  PIN E2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 40.600 110.000 41.160 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 42.840 110.000 43.400 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 46.200 110.000 46.760 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 49.560 110.000 50.120 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 52.920 110.000 53.480 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 55.160 110.000 55.720 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 58.520 110.000 59.080 ;
    END
  END E2BEGb[7]
  PIN E6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 110.040 110.000 110.600 ;
    END
  END E6BEG[0]
  PIN E6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 140.280 110.000 140.840 ;
    END
  END E6BEG[10]
  PIN E6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 143.640 110.000 144.200 ;
    END
  END E6BEG[11]
  PIN E6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 113.400 110.000 113.960 ;
    END
  END E6BEG[1]
  PIN E6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 116.760 110.000 117.320 ;
    END
  END E6BEG[2]
  PIN E6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 119.000 110.000 119.560 ;
    END
  END E6BEG[3]
  PIN E6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 122.360 110.000 122.920 ;
    END
  END E6BEG[4]
  PIN E6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 125.720 110.000 126.280 ;
    END
  END E6BEG[5]
  PIN E6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 127.960 110.000 128.520 ;
    END
  END E6BEG[6]
  PIN E6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 131.320 110.000 131.880 ;
    END
  END E6BEG[7]
  PIN E6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 134.680 110.000 135.240 ;
    END
  END E6BEG[8]
  PIN E6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 136.920 110.000 137.480 ;
    END
  END E6BEG[9]
  PIN EE4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 61.880 110.000 62.440 ;
    END
  END EE4BEG[0]
  PIN EE4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 92.120 110.000 92.680 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 95.480 110.000 96.040 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 97.720 110.000 98.280 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 101.080 110.000 101.640 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 104.440 110.000 105.000 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 106.680 110.000 107.240 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 64.120 110.000 64.680 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 67.480 110.000 68.040 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 70.840 110.000 71.400 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 74.200 110.000 74.760 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 76.440 110.000 77.000 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 79.800 110.000 80.360 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 83.160 110.000 83.720 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 85.400 110.000 85.960 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 88.760 110.000 89.320 ;
    END
  END EE4BEG[9]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 119.000 2.000 119.560 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 204.120 2.000 204.680 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 211.960 2.000 212.520 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 220.920 2.000 221.480 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 228.760 2.000 229.320 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 237.720 2.000 238.280 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 245.560 2.000 246.120 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 254.520 2.000 255.080 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.360 2.000 262.920 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 271.320 2.000 271.880 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 279.160 2.000 279.720 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.960 2.000 128.520 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 288.120 2.000 288.680 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 297.080 2.000 297.640 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 304.920 2.000 305.480 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 313.880 2.000 314.440 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 321.720 2.000 322.280 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 330.680 2.000 331.240 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 338.520 2.000 339.080 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 347.480 2.000 348.040 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 355.320 2.000 355.880 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 364.280 2.000 364.840 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 135.800 2.000 136.360 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 372.120 2.000 372.680 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 381.080 2.000 381.640 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 144.760 2.000 145.320 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 152.600 2.000 153.160 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 161.560 2.000 162.120 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 169.400 2.000 169.960 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 178.360 2.000 178.920 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 186.200 2.000 186.760 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 195.160 2.000 195.720 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 292.600 110.000 293.160 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 322.840 110.000 323.400 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 326.200 110.000 326.760 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 328.440 110.000 329.000 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 331.800 110.000 332.360 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 335.160 110.000 335.720 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 337.400 110.000 337.960 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 340.760 110.000 341.320 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 344.120 110.000 344.680 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 347.480 110.000 348.040 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 349.720 110.000 350.280 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 294.840 110.000 295.400 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 353.080 110.000 353.640 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 356.440 110.000 357.000 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 358.680 110.000 359.240 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 362.040 110.000 362.600 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 365.400 110.000 365.960 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 368.760 110.000 369.320 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 371.000 110.000 371.560 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 374.360 110.000 374.920 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 377.720 110.000 378.280 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 379.960 110.000 380.520 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 298.200 110.000 298.760 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 383.320 110.000 383.880 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 386.680 110.000 387.240 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 301.560 110.000 302.120 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 304.920 110.000 305.480 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 307.160 110.000 307.720 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 310.520 110.000 311.080 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 313.880 110.000 314.440 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 316.120 110.000 316.680 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 319.480 110.000 320.040 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 5.880 0.000 6.440 2.000 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.400 0.000 57.960 2.000 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.000 0.000 63.560 2.000 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 68.600 0.000 69.160 2.000 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.080 0.000 73.640 2.000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 78.680 0.000 79.240 2.000 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 83.160 0.000 83.720 2.000 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 88.760 0.000 89.320 2.000 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.360 0.000 94.920 2.000 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 98.840 0.000 99.400 2.000 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.440 0.000 105.000 2.000 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 11.480 0.000 12.040 2.000 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 15.960 0.000 16.520 2.000 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 21.560 0.000 22.120 2.000 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 27.160 0.000 27.720 2.000 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 31.640 0.000 32.200 2.000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 37.240 0.000 37.800 2.000 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.720 0.000 42.280 2.000 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.320 0.000 47.880 2.000 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 52.920 0.000 53.480 2.000 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 5.880 388.000 6.440 390.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.400 388.000 57.960 390.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.000 388.000 63.560 390.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 68.600 388.000 69.160 390.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.080 388.000 73.640 390.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 78.680 388.000 79.240 390.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 83.160 388.000 83.720 390.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 88.760 388.000 89.320 390.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.360 388.000 94.920 390.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 98.840 388.000 99.400 390.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.440 388.000 105.000 390.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 11.480 388.000 12.040 390.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 15.960 388.000 16.520 390.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 21.560 388.000 22.120 390.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 27.160 388.000 27.720 390.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 31.640 388.000 32.200 390.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 37.240 388.000 37.800 390.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.720 388.000 42.280 390.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.320 388.000 47.880 390.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 52.920 388.000 53.480 390.000 ;
    END
  END FrameStrobe_O[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1.400 0.000 1.960 2.000 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1.400 388.000 1.960 390.000 ;
    END
  END UserCLKo
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 17.960 7.540 19.560 380.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 42.040 7.540 43.640 380.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 66.120 7.540 67.720 380.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 90.200 7.540 91.800 380.540 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 30.000 7.540 31.600 380.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 54.080 7.540 55.680 380.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 78.160 7.540 79.760 380.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 102.240 7.540 103.840 380.540 ;
    END
  END VSS
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 147.000 110.000 147.560 ;
    END
  END W1END[0]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 149.240 110.000 149.800 ;
    END
  END W1END[1]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 152.600 110.000 153.160 ;
    END
  END W1END[2]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 155.960 110.000 156.520 ;
    END
  END W1END[3]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 182.840 110.000 183.400 ;
    END
  END W2END[0]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 186.200 110.000 186.760 ;
    END
  END W2END[1]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 189.560 110.000 190.120 ;
    END
  END W2END[2]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 191.800 110.000 192.360 ;
    END
  END W2END[3]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 195.160 110.000 195.720 ;
    END
  END W2END[4]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 198.520 110.000 199.080 ;
    END
  END W2END[5]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 200.760 110.000 201.320 ;
    END
  END W2END[6]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 204.120 110.000 204.680 ;
    END
  END W2END[7]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 158.200 110.000 158.760 ;
    END
  END W2MID[0]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 161.560 110.000 162.120 ;
    END
  END W2MID[1]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 164.920 110.000 165.480 ;
    END
  END W2MID[2]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 168.280 110.000 168.840 ;
    END
  END W2MID[3]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 170.520 110.000 171.080 ;
    END
  END W2MID[4]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 173.880 110.000 174.440 ;
    END
  END W2MID[5]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 177.240 110.000 177.800 ;
    END
  END W2MID[6]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 179.480 110.000 180.040 ;
    END
  END W2MID[7]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 255.640 110.000 256.200 ;
    END
  END W6END[0]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 285.880 110.000 286.440 ;
    END
  END W6END[10]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 289.240 110.000 289.800 ;
    END
  END W6END[11]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 259.000 110.000 259.560 ;
    END
  END W6END[1]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 262.360 110.000 262.920 ;
    END
  END W6END[2]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 264.600 110.000 265.160 ;
    END
  END W6END[3]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 267.960 110.000 268.520 ;
    END
  END W6END[4]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 271.320 110.000 271.880 ;
    END
  END W6END[5]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 273.560 110.000 274.120 ;
    END
  END W6END[6]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 276.920 110.000 277.480 ;
    END
  END W6END[7]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 280.280 110.000 280.840 ;
    END
  END W6END[8]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 283.640 110.000 284.200 ;
    END
  END W6END[9]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 207.480 110.000 208.040 ;
    END
  END WW4END[0]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 237.720 110.000 238.280 ;
    END
  END WW4END[10]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 241.080 110.000 241.640 ;
    END
  END WW4END[11]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 243.320 110.000 243.880 ;
    END
  END WW4END[12]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 246.680 110.000 247.240 ;
    END
  END WW4END[13]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 250.040 110.000 250.600 ;
    END
  END WW4END[14]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 253.400 110.000 253.960 ;
    END
  END WW4END[15]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 210.840 110.000 211.400 ;
    END
  END WW4END[1]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 213.080 110.000 213.640 ;
    END
  END WW4END[2]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 216.440 110.000 217.000 ;
    END
  END WW4END[3]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 219.800 110.000 220.360 ;
    END
  END WW4END[4]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 222.040 110.000 222.600 ;
    END
  END WW4END[5]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 225.400 110.000 225.960 ;
    END
  END WW4END[6]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 228.760 110.000 229.320 ;
    END
  END WW4END[7]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 232.120 110.000 232.680 ;
    END
  END WW4END[8]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 234.360 110.000 234.920 ;
    END
  END WW4END[9]
  OBS
      LAYER Metal1 ;
        RECT 6.720 4.070 109.670 381.210 ;
      LAYER Metal2 ;
        RECT 0.140 387.700 1.100 388.500 ;
        RECT 2.260 387.700 5.580 388.500 ;
        RECT 6.740 387.700 11.180 388.500 ;
        RECT 12.340 387.700 15.660 388.500 ;
        RECT 16.820 387.700 21.260 388.500 ;
        RECT 22.420 387.700 26.860 388.500 ;
        RECT 28.020 387.700 31.340 388.500 ;
        RECT 32.500 387.700 36.940 388.500 ;
        RECT 38.100 387.700 41.420 388.500 ;
        RECT 42.580 387.700 47.020 388.500 ;
        RECT 48.180 387.700 52.620 388.500 ;
        RECT 53.780 387.700 57.100 388.500 ;
        RECT 58.260 387.700 62.700 388.500 ;
        RECT 63.860 387.700 68.300 388.500 ;
        RECT 69.460 387.700 72.780 388.500 ;
        RECT 73.940 387.700 78.380 388.500 ;
        RECT 79.540 387.700 82.860 388.500 ;
        RECT 84.020 387.700 88.460 388.500 ;
        RECT 89.620 387.700 94.060 388.500 ;
        RECT 95.220 387.700 98.540 388.500 ;
        RECT 99.700 387.700 104.140 388.500 ;
        RECT 105.300 387.700 109.620 388.500 ;
        RECT 0.140 2.300 109.620 387.700 ;
        RECT 0.140 1.260 1.100 2.300 ;
        RECT 2.260 1.260 5.580 2.300 ;
        RECT 6.740 1.260 11.180 2.300 ;
        RECT 12.340 1.260 15.660 2.300 ;
        RECT 16.820 1.260 21.260 2.300 ;
        RECT 22.420 1.260 26.860 2.300 ;
        RECT 28.020 1.260 31.340 2.300 ;
        RECT 32.500 1.260 36.940 2.300 ;
        RECT 38.100 1.260 41.420 2.300 ;
        RECT 42.580 1.260 47.020 2.300 ;
        RECT 48.180 1.260 52.620 2.300 ;
        RECT 53.780 1.260 57.100 2.300 ;
        RECT 58.260 1.260 62.700 2.300 ;
        RECT 63.860 1.260 68.300 2.300 ;
        RECT 69.460 1.260 72.780 2.300 ;
        RECT 73.940 1.260 78.380 2.300 ;
        RECT 79.540 1.260 82.860 2.300 ;
        RECT 84.020 1.260 88.460 2.300 ;
        RECT 89.620 1.260 94.060 2.300 ;
        RECT 95.220 1.260 98.540 2.300 ;
        RECT 99.700 1.260 104.140 2.300 ;
        RECT 105.300 1.260 109.620 2.300 ;
      LAYER Metal3 ;
        RECT 0.090 386.380 107.700 386.820 ;
        RECT 0.090 384.180 109.670 386.380 ;
        RECT 0.090 383.020 107.700 384.180 ;
        RECT 0.090 381.940 109.670 383.020 ;
        RECT 2.300 380.820 109.670 381.940 ;
        RECT 2.300 380.780 107.700 380.820 ;
        RECT 0.090 379.660 107.700 380.780 ;
        RECT 0.090 378.580 109.670 379.660 ;
        RECT 0.090 377.420 107.700 378.580 ;
        RECT 0.090 375.220 109.670 377.420 ;
        RECT 0.090 374.060 107.700 375.220 ;
        RECT 0.090 372.980 109.670 374.060 ;
        RECT 2.300 371.860 109.670 372.980 ;
        RECT 2.300 371.820 107.700 371.860 ;
        RECT 0.090 370.700 107.700 371.820 ;
        RECT 0.090 369.620 109.670 370.700 ;
        RECT 0.090 368.460 107.700 369.620 ;
        RECT 0.090 366.260 109.670 368.460 ;
        RECT 0.090 365.140 107.700 366.260 ;
        RECT 2.300 365.100 107.700 365.140 ;
        RECT 2.300 363.980 109.670 365.100 ;
        RECT 0.090 362.900 109.670 363.980 ;
        RECT 0.090 361.740 107.700 362.900 ;
        RECT 0.090 359.540 109.670 361.740 ;
        RECT 0.090 358.380 107.700 359.540 ;
        RECT 0.090 357.300 109.670 358.380 ;
        RECT 0.090 356.180 107.700 357.300 ;
        RECT 2.300 356.140 107.700 356.180 ;
        RECT 2.300 355.020 109.670 356.140 ;
        RECT 0.090 353.940 109.670 355.020 ;
        RECT 0.090 352.780 107.700 353.940 ;
        RECT 0.090 350.580 109.670 352.780 ;
        RECT 0.090 349.420 107.700 350.580 ;
        RECT 0.090 348.340 109.670 349.420 ;
        RECT 2.300 347.180 107.700 348.340 ;
        RECT 0.090 344.980 109.670 347.180 ;
        RECT 0.090 343.820 107.700 344.980 ;
        RECT 0.090 341.620 109.670 343.820 ;
        RECT 0.090 340.460 107.700 341.620 ;
        RECT 0.090 339.380 109.670 340.460 ;
        RECT 2.300 338.260 109.670 339.380 ;
        RECT 2.300 338.220 107.700 338.260 ;
        RECT 0.090 337.100 107.700 338.220 ;
        RECT 0.090 336.020 109.670 337.100 ;
        RECT 0.090 334.860 107.700 336.020 ;
        RECT 0.090 332.660 109.670 334.860 ;
        RECT 0.090 331.540 107.700 332.660 ;
        RECT 2.300 331.500 107.700 331.540 ;
        RECT 2.300 330.380 109.670 331.500 ;
        RECT 0.090 329.300 109.670 330.380 ;
        RECT 0.090 328.140 107.700 329.300 ;
        RECT 0.090 327.060 109.670 328.140 ;
        RECT 0.090 325.900 107.700 327.060 ;
        RECT 0.090 323.700 109.670 325.900 ;
        RECT 0.090 322.580 107.700 323.700 ;
        RECT 2.300 322.540 107.700 322.580 ;
        RECT 2.300 321.420 109.670 322.540 ;
        RECT 0.090 320.340 109.670 321.420 ;
        RECT 0.090 319.180 107.700 320.340 ;
        RECT 0.090 316.980 109.670 319.180 ;
        RECT 0.090 315.820 107.700 316.980 ;
        RECT 0.090 314.740 109.670 315.820 ;
        RECT 2.300 313.580 107.700 314.740 ;
        RECT 0.090 311.380 109.670 313.580 ;
        RECT 0.090 310.220 107.700 311.380 ;
        RECT 0.090 308.020 109.670 310.220 ;
        RECT 0.090 306.860 107.700 308.020 ;
        RECT 0.090 305.780 109.670 306.860 ;
        RECT 2.300 304.620 107.700 305.780 ;
        RECT 0.090 302.420 109.670 304.620 ;
        RECT 0.090 301.260 107.700 302.420 ;
        RECT 0.090 299.060 109.670 301.260 ;
        RECT 0.090 297.940 107.700 299.060 ;
        RECT 2.300 297.900 107.700 297.940 ;
        RECT 2.300 296.780 109.670 297.900 ;
        RECT 0.090 295.700 109.670 296.780 ;
        RECT 0.090 294.540 107.700 295.700 ;
        RECT 0.090 293.460 109.670 294.540 ;
        RECT 0.090 292.300 107.700 293.460 ;
        RECT 0.090 290.100 109.670 292.300 ;
        RECT 0.090 288.980 107.700 290.100 ;
        RECT 2.300 288.940 107.700 288.980 ;
        RECT 2.300 287.820 109.670 288.940 ;
        RECT 0.090 286.740 109.670 287.820 ;
        RECT 0.090 285.580 107.700 286.740 ;
        RECT 0.090 284.500 109.670 285.580 ;
        RECT 0.090 283.340 107.700 284.500 ;
        RECT 0.090 281.140 109.670 283.340 ;
        RECT 0.090 280.020 107.700 281.140 ;
        RECT 2.300 279.980 107.700 280.020 ;
        RECT 2.300 278.860 109.670 279.980 ;
        RECT 0.090 277.780 109.670 278.860 ;
        RECT 0.090 276.620 107.700 277.780 ;
        RECT 0.090 274.420 109.670 276.620 ;
        RECT 0.090 273.260 107.700 274.420 ;
        RECT 0.090 272.180 109.670 273.260 ;
        RECT 2.300 271.020 107.700 272.180 ;
        RECT 0.090 268.820 109.670 271.020 ;
        RECT 0.090 267.660 107.700 268.820 ;
        RECT 0.090 265.460 109.670 267.660 ;
        RECT 0.090 264.300 107.700 265.460 ;
        RECT 0.090 263.220 109.670 264.300 ;
        RECT 2.300 262.060 107.700 263.220 ;
        RECT 0.090 259.860 109.670 262.060 ;
        RECT 0.090 258.700 107.700 259.860 ;
        RECT 0.090 256.500 109.670 258.700 ;
        RECT 0.090 255.380 107.700 256.500 ;
        RECT 2.300 255.340 107.700 255.380 ;
        RECT 2.300 254.260 109.670 255.340 ;
        RECT 2.300 254.220 107.700 254.260 ;
        RECT 0.090 253.100 107.700 254.220 ;
        RECT 0.090 250.900 109.670 253.100 ;
        RECT 0.090 249.740 107.700 250.900 ;
        RECT 0.090 247.540 109.670 249.740 ;
        RECT 0.090 246.420 107.700 247.540 ;
        RECT 2.300 246.380 107.700 246.420 ;
        RECT 2.300 245.260 109.670 246.380 ;
        RECT 0.090 244.180 109.670 245.260 ;
        RECT 0.090 243.020 107.700 244.180 ;
        RECT 0.090 241.940 109.670 243.020 ;
        RECT 0.090 240.780 107.700 241.940 ;
        RECT 0.090 238.580 109.670 240.780 ;
        RECT 2.300 237.420 107.700 238.580 ;
        RECT 0.090 235.220 109.670 237.420 ;
        RECT 0.090 234.060 107.700 235.220 ;
        RECT 0.090 232.980 109.670 234.060 ;
        RECT 0.090 231.820 107.700 232.980 ;
        RECT 0.090 229.620 109.670 231.820 ;
        RECT 2.300 228.460 107.700 229.620 ;
        RECT 0.090 226.260 109.670 228.460 ;
        RECT 0.090 225.100 107.700 226.260 ;
        RECT 0.090 222.900 109.670 225.100 ;
        RECT 0.090 221.780 107.700 222.900 ;
        RECT 2.300 221.740 107.700 221.780 ;
        RECT 2.300 220.660 109.670 221.740 ;
        RECT 2.300 220.620 107.700 220.660 ;
        RECT 0.090 219.500 107.700 220.620 ;
        RECT 0.090 217.300 109.670 219.500 ;
        RECT 0.090 216.140 107.700 217.300 ;
        RECT 0.090 213.940 109.670 216.140 ;
        RECT 0.090 212.820 107.700 213.940 ;
        RECT 2.300 212.780 107.700 212.820 ;
        RECT 2.300 211.700 109.670 212.780 ;
        RECT 2.300 211.660 107.700 211.700 ;
        RECT 0.090 210.540 107.700 211.660 ;
        RECT 0.090 208.340 109.670 210.540 ;
        RECT 0.090 207.180 107.700 208.340 ;
        RECT 0.090 204.980 109.670 207.180 ;
        RECT 2.300 203.820 107.700 204.980 ;
        RECT 0.090 201.620 109.670 203.820 ;
        RECT 0.090 200.460 107.700 201.620 ;
        RECT 0.090 199.380 109.670 200.460 ;
        RECT 0.090 198.220 107.700 199.380 ;
        RECT 0.090 196.020 109.670 198.220 ;
        RECT 2.300 194.860 107.700 196.020 ;
        RECT 0.090 192.660 109.670 194.860 ;
        RECT 0.090 191.500 107.700 192.660 ;
        RECT 0.090 190.420 109.670 191.500 ;
        RECT 0.090 189.260 107.700 190.420 ;
        RECT 0.090 187.060 109.670 189.260 ;
        RECT 2.300 185.900 107.700 187.060 ;
        RECT 0.090 183.700 109.670 185.900 ;
        RECT 0.090 182.540 107.700 183.700 ;
        RECT 0.090 180.340 109.670 182.540 ;
        RECT 0.090 179.220 107.700 180.340 ;
        RECT 2.300 179.180 107.700 179.220 ;
        RECT 2.300 178.100 109.670 179.180 ;
        RECT 2.300 178.060 107.700 178.100 ;
        RECT 0.090 176.940 107.700 178.060 ;
        RECT 0.090 174.740 109.670 176.940 ;
        RECT 0.090 173.580 107.700 174.740 ;
        RECT 0.090 171.380 109.670 173.580 ;
        RECT 0.090 170.260 107.700 171.380 ;
        RECT 2.300 170.220 107.700 170.260 ;
        RECT 2.300 169.140 109.670 170.220 ;
        RECT 2.300 169.100 107.700 169.140 ;
        RECT 0.090 167.980 107.700 169.100 ;
        RECT 0.090 165.780 109.670 167.980 ;
        RECT 0.090 164.620 107.700 165.780 ;
        RECT 0.090 162.420 109.670 164.620 ;
        RECT 2.300 161.260 107.700 162.420 ;
        RECT 0.090 159.060 109.670 161.260 ;
        RECT 0.090 157.900 107.700 159.060 ;
        RECT 0.090 156.820 109.670 157.900 ;
        RECT 0.090 155.660 107.700 156.820 ;
        RECT 0.090 153.460 109.670 155.660 ;
        RECT 2.300 152.300 107.700 153.460 ;
        RECT 0.090 150.100 109.670 152.300 ;
        RECT 0.090 148.940 107.700 150.100 ;
        RECT 0.090 147.860 109.670 148.940 ;
        RECT 0.090 146.700 107.700 147.860 ;
        RECT 0.090 145.620 109.670 146.700 ;
        RECT 2.300 144.500 109.670 145.620 ;
        RECT 2.300 144.460 107.700 144.500 ;
        RECT 0.090 143.340 107.700 144.460 ;
        RECT 0.090 141.140 109.670 143.340 ;
        RECT 0.090 139.980 107.700 141.140 ;
        RECT 0.090 137.780 109.670 139.980 ;
        RECT 0.090 136.660 107.700 137.780 ;
        RECT 2.300 136.620 107.700 136.660 ;
        RECT 2.300 135.540 109.670 136.620 ;
        RECT 2.300 135.500 107.700 135.540 ;
        RECT 0.090 134.380 107.700 135.500 ;
        RECT 0.090 132.180 109.670 134.380 ;
        RECT 0.090 131.020 107.700 132.180 ;
        RECT 0.090 128.820 109.670 131.020 ;
        RECT 2.300 127.660 107.700 128.820 ;
        RECT 0.090 126.580 109.670 127.660 ;
        RECT 0.090 125.420 107.700 126.580 ;
        RECT 0.090 123.220 109.670 125.420 ;
        RECT 0.090 122.060 107.700 123.220 ;
        RECT 0.090 119.860 109.670 122.060 ;
        RECT 2.300 118.700 107.700 119.860 ;
        RECT 0.090 117.620 109.670 118.700 ;
        RECT 0.090 116.460 107.700 117.620 ;
        RECT 0.090 114.260 109.670 116.460 ;
        RECT 0.090 113.100 107.700 114.260 ;
        RECT 0.090 112.020 109.670 113.100 ;
        RECT 2.300 110.900 109.670 112.020 ;
        RECT 2.300 110.860 107.700 110.900 ;
        RECT 0.090 109.740 107.700 110.860 ;
        RECT 0.090 107.540 109.670 109.740 ;
        RECT 0.090 106.380 107.700 107.540 ;
        RECT 0.090 105.300 109.670 106.380 ;
        RECT 0.090 104.140 107.700 105.300 ;
        RECT 0.090 103.060 109.670 104.140 ;
        RECT 2.300 101.940 109.670 103.060 ;
        RECT 2.300 101.900 107.700 101.940 ;
        RECT 0.090 100.780 107.700 101.900 ;
        RECT 0.090 98.580 109.670 100.780 ;
        RECT 0.090 97.420 107.700 98.580 ;
        RECT 0.090 96.340 109.670 97.420 ;
        RECT 0.090 95.180 107.700 96.340 ;
        RECT 0.090 94.100 109.670 95.180 ;
        RECT 2.300 92.980 109.670 94.100 ;
        RECT 2.300 92.940 107.700 92.980 ;
        RECT 0.090 91.820 107.700 92.940 ;
        RECT 0.090 89.620 109.670 91.820 ;
        RECT 0.090 88.460 107.700 89.620 ;
        RECT 0.090 86.260 109.670 88.460 ;
        RECT 2.300 85.100 107.700 86.260 ;
        RECT 0.090 84.020 109.670 85.100 ;
        RECT 0.090 82.860 107.700 84.020 ;
        RECT 0.090 80.660 109.670 82.860 ;
        RECT 0.090 79.500 107.700 80.660 ;
        RECT 0.090 77.300 109.670 79.500 ;
        RECT 2.300 76.140 107.700 77.300 ;
        RECT 0.090 75.060 109.670 76.140 ;
        RECT 0.090 73.900 107.700 75.060 ;
        RECT 0.090 71.700 109.670 73.900 ;
        RECT 0.090 70.540 107.700 71.700 ;
        RECT 0.090 69.460 109.670 70.540 ;
        RECT 2.300 68.340 109.670 69.460 ;
        RECT 2.300 68.300 107.700 68.340 ;
        RECT 0.090 67.180 107.700 68.300 ;
        RECT 0.090 64.980 109.670 67.180 ;
        RECT 0.090 63.820 107.700 64.980 ;
        RECT 0.090 62.740 109.670 63.820 ;
        RECT 0.090 61.580 107.700 62.740 ;
        RECT 0.090 60.500 109.670 61.580 ;
        RECT 2.300 59.380 109.670 60.500 ;
        RECT 2.300 59.340 107.700 59.380 ;
        RECT 0.090 58.220 107.700 59.340 ;
        RECT 0.090 56.020 109.670 58.220 ;
        RECT 0.090 54.860 107.700 56.020 ;
        RECT 0.090 53.780 109.670 54.860 ;
        RECT 0.090 52.660 107.700 53.780 ;
        RECT 2.300 52.620 107.700 52.660 ;
        RECT 2.300 51.500 109.670 52.620 ;
        RECT 0.090 50.420 109.670 51.500 ;
        RECT 0.090 49.260 107.700 50.420 ;
        RECT 0.090 47.060 109.670 49.260 ;
        RECT 0.090 45.900 107.700 47.060 ;
        RECT 0.090 43.700 109.670 45.900 ;
        RECT 2.300 42.540 107.700 43.700 ;
        RECT 0.090 41.460 109.670 42.540 ;
        RECT 0.090 40.300 107.700 41.460 ;
        RECT 0.090 38.100 109.670 40.300 ;
        RECT 0.090 36.940 107.700 38.100 ;
        RECT 0.090 35.860 109.670 36.940 ;
        RECT 2.300 34.740 109.670 35.860 ;
        RECT 2.300 34.700 107.700 34.740 ;
        RECT 0.090 33.580 107.700 34.700 ;
        RECT 0.090 32.500 109.670 33.580 ;
        RECT 0.090 31.340 107.700 32.500 ;
        RECT 0.090 29.140 109.670 31.340 ;
        RECT 0.090 27.980 107.700 29.140 ;
        RECT 0.090 26.900 109.670 27.980 ;
        RECT 2.300 25.780 109.670 26.900 ;
        RECT 2.300 25.740 107.700 25.780 ;
        RECT 0.090 24.620 107.700 25.740 ;
        RECT 0.090 22.420 109.670 24.620 ;
        RECT 0.090 21.260 107.700 22.420 ;
        RECT 0.090 20.180 109.670 21.260 ;
        RECT 0.090 19.060 107.700 20.180 ;
        RECT 2.300 19.020 107.700 19.060 ;
        RECT 2.300 17.900 109.670 19.020 ;
        RECT 0.090 16.820 109.670 17.900 ;
        RECT 0.090 15.660 107.700 16.820 ;
        RECT 0.090 13.460 109.670 15.660 ;
        RECT 0.090 12.300 107.700 13.460 ;
        RECT 0.090 11.220 109.670 12.300 ;
        RECT 0.090 10.100 107.700 11.220 ;
        RECT 2.300 10.060 107.700 10.100 ;
        RECT 2.300 8.940 109.670 10.060 ;
        RECT 0.090 7.860 109.670 8.940 ;
        RECT 0.090 6.700 107.700 7.860 ;
        RECT 0.090 4.500 109.670 6.700 ;
        RECT 0.090 3.340 107.700 4.500 ;
        RECT 0.090 2.260 109.670 3.340 ;
        RECT 2.300 1.820 107.700 2.260 ;
      LAYER Metal4 ;
        RECT 24.220 7.240 29.700 376.230 ;
        RECT 31.900 7.240 41.740 376.230 ;
        RECT 43.940 7.240 53.780 376.230 ;
        RECT 55.980 7.240 65.820 376.230 ;
        RECT 68.020 7.240 77.860 376.230 ;
        RECT 80.060 7.240 89.900 376.230 ;
        RECT 92.100 7.240 101.940 376.230 ;
        RECT 104.140 7.240 107.380 376.230 ;
        RECT 24.220 2.890 107.380 7.240 ;
  END
END W_IO
END LIBRARY

