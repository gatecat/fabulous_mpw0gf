VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO S_term_single2
  CLASS BLOCK ;
  FOREIGN S_term_single2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 450.000 BY 180.000 ;
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 22.680 0.000 23.240 2.000 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 235.480 0.000 236.040 2.000 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 256.760 0.000 257.320 2.000 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.040 0.000 278.600 2.000 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 299.320 0.000 299.880 2.000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 320.600 0.000 321.160 2.000 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 341.880 0.000 342.440 2.000 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 363.160 0.000 363.720 2.000 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 384.440 0.000 385.000 2.000 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 405.720 0.000 406.280 2.000 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 427.000 0.000 427.560 2.000 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.960 0.000 44.520 2.000 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 65.240 0.000 65.800 2.000 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 86.520 0.000 87.080 2.000 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.800 0.000 108.360 2.000 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 129.080 0.000 129.640 2.000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 150.360 0.000 150.920 2.000 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.640 0.000 172.200 2.000 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 192.920 0.000 193.480 2.000 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 214.200 0.000 214.760 2.000 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 377.720 178.000 378.280 180.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 413.560 178.000 414.120 180.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 416.920 178.000 417.480 180.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 420.280 178.000 420.840 180.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 423.640 178.000 424.200 180.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 427.000 178.000 427.560 180.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 431.480 178.000 432.040 180.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 434.840 178.000 435.400 180.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 438.200 178.000 438.760 180.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 441.560 178.000 442.120 180.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 444.920 178.000 445.480 180.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 381.080 178.000 381.640 180.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 384.440 178.000 385.000 180.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 387.800 178.000 388.360 180.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 391.160 178.000 391.720 180.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 395.640 178.000 396.200 180.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 399.000 178.000 399.560 180.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 402.360 178.000 402.920 180.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 405.720 178.000 406.280 180.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 409.080 178.000 409.640 180.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1.400 178.000 1.960 180.000 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 4.760 178.000 5.320 180.000 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 8.120 178.000 8.680 180.000 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 11.480 178.000 12.040 180.000 ;
    END
  END N1BEG[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 14.840 178.000 15.400 180.000 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 19.320 178.000 19.880 180.000 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 22.680 178.000 23.240 180.000 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.040 178.000 26.600 180.000 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 29.400 178.000 29.960 180.000 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 32.760 178.000 33.320 180.000 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 37.240 178.000 37.800 180.000 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.600 178.000 41.160 180.000 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.960 178.000 44.520 180.000 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.320 178.000 47.880 180.000 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.680 178.000 51.240 180.000 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 55.160 178.000 55.720 180.000 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 58.520 178.000 59.080 180.000 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 61.880 178.000 62.440 180.000 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 65.240 178.000 65.800 180.000 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 68.600 178.000 69.160 180.000 ;
    END
  END N2BEGb[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.080 178.000 73.640 180.000 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 108.920 178.000 109.480 180.000 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 112.280 178.000 112.840 180.000 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 115.640 178.000 116.200 180.000 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 119.000 178.000 119.560 180.000 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 122.360 178.000 122.920 180.000 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 126.840 178.000 127.400 180.000 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 76.440 178.000 77.000 180.000 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 79.800 178.000 80.360 180.000 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 83.160 178.000 83.720 180.000 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 86.520 178.000 87.080 180.000 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 91.000 178.000 91.560 180.000 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.360 178.000 94.920 180.000 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.720 178.000 98.280 180.000 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 101.080 178.000 101.640 180.000 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.440 178.000 105.000 180.000 ;
    END
  END N4BEG[9]
  PIN NN4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 130.200 178.000 130.760 180.000 ;
    END
  END NN4BEG[0]
  PIN NN4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 166.040 178.000 166.600 180.000 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 169.400 178.000 169.960 180.000 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 172.760 178.000 173.320 180.000 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 176.120 178.000 176.680 180.000 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 180.600 178.000 181.160 180.000 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 183.960 178.000 184.520 180.000 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 133.560 178.000 134.120 180.000 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 136.920 178.000 137.480 180.000 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 140.280 178.000 140.840 180.000 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.760 178.000 145.320 180.000 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 148.120 178.000 148.680 180.000 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.480 178.000 152.040 180.000 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.840 178.000 155.400 180.000 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 158.200 178.000 158.760 180.000 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 162.680 178.000 163.240 180.000 ;
    END
  END NN4BEG[9]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 187.320 178.000 187.880 180.000 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 190.680 178.000 191.240 180.000 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.040 178.000 194.600 180.000 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 198.520 178.000 199.080 180.000 ;
    END
  END S1END[3]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 229.880 178.000 230.440 180.000 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.360 178.000 234.920 180.000 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 237.720 178.000 238.280 180.000 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.080 178.000 241.640 180.000 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 244.440 178.000 245.000 180.000 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 247.800 178.000 248.360 180.000 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 252.280 178.000 252.840 180.000 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 255.640 178.000 256.200 180.000 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.880 178.000 202.440 180.000 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 205.240 178.000 205.800 180.000 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 208.600 178.000 209.160 180.000 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.960 178.000 212.520 180.000 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 216.440 178.000 217.000 180.000 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 219.800 178.000 220.360 180.000 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 223.160 178.000 223.720 180.000 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 226.520 178.000 227.080 180.000 ;
    END
  END S2MID[7]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 259.000 178.000 259.560 180.000 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 294.840 178.000 295.400 180.000 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 298.200 178.000 298.760 180.000 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 301.560 178.000 302.120 180.000 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 306.040 178.000 306.600 180.000 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 309.400 178.000 309.960 180.000 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 312.760 178.000 313.320 180.000 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.360 178.000 262.920 180.000 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 265.720 178.000 266.280 180.000 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 270.200 178.000 270.760 180.000 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 273.560 178.000 274.120 180.000 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 276.920 178.000 277.480 180.000 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 280.280 178.000 280.840 180.000 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 283.640 178.000 284.200 180.000 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.120 178.000 288.680 180.000 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 291.480 178.000 292.040 180.000 ;
    END
  END S4END[9]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 316.120 178.000 316.680 180.000 ;
    END
  END SS4END[0]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 351.960 178.000 352.520 180.000 ;
    END
  END SS4END[10]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 355.320 178.000 355.880 180.000 ;
    END
  END SS4END[11]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 359.800 178.000 360.360 180.000 ;
    END
  END SS4END[12]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 363.160 178.000 363.720 180.000 ;
    END
  END SS4END[13]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 366.520 178.000 367.080 180.000 ;
    END
  END SS4END[14]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 369.880 178.000 370.440 180.000 ;
    END
  END SS4END[15]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 319.480 178.000 320.040 180.000 ;
    END
  END SS4END[1]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 323.960 178.000 324.520 180.000 ;
    END
  END SS4END[2]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 327.320 178.000 327.880 180.000 ;
    END
  END SS4END[3]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 330.680 178.000 331.240 180.000 ;
    END
  END SS4END[4]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 334.040 178.000 334.600 180.000 ;
    END
  END SS4END[5]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 337.400 178.000 337.960 180.000 ;
    END
  END SS4END[6]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 341.880 178.000 342.440 180.000 ;
    END
  END SS4END[7]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 345.240 178.000 345.800 180.000 ;
    END
  END SS4END[8]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 348.600 178.000 349.160 180.000 ;
    END
  END SS4END[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1.400 0.000 1.960 2.000 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 373.240 178.000 373.800 180.000 ;
    END
  END UserCLKo
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 60.445 7.540 62.045 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 169.500 7.540 171.100 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 278.555 7.540 280.155 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 387.610 7.540 389.210 168.860 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 114.970 7.540 116.570 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 224.025 7.540 225.625 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 333.080 7.540 334.680 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 442.135 7.540 443.735 168.860 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 7.540 443.735 172.890 ;
      LAYER Metal2 ;
        RECT 2.260 177.700 4.460 179.110 ;
        RECT 5.620 177.700 7.820 179.110 ;
        RECT 8.980 177.700 11.180 179.110 ;
        RECT 12.340 177.700 14.540 179.110 ;
        RECT 15.700 177.700 19.020 179.110 ;
        RECT 20.180 177.700 22.380 179.110 ;
        RECT 23.540 177.700 25.740 179.110 ;
        RECT 26.900 177.700 29.100 179.110 ;
        RECT 30.260 177.700 32.460 179.110 ;
        RECT 33.620 177.700 36.940 179.110 ;
        RECT 38.100 177.700 40.300 179.110 ;
        RECT 41.460 177.700 43.660 179.110 ;
        RECT 44.820 177.700 47.020 179.110 ;
        RECT 48.180 177.700 50.380 179.110 ;
        RECT 51.540 177.700 54.860 179.110 ;
        RECT 56.020 177.700 58.220 179.110 ;
        RECT 59.380 177.700 61.580 179.110 ;
        RECT 62.740 177.700 64.940 179.110 ;
        RECT 66.100 177.700 68.300 179.110 ;
        RECT 69.460 177.700 72.780 179.110 ;
        RECT 73.940 177.700 76.140 179.110 ;
        RECT 77.300 177.700 79.500 179.110 ;
        RECT 80.660 177.700 82.860 179.110 ;
        RECT 84.020 177.700 86.220 179.110 ;
        RECT 87.380 177.700 90.700 179.110 ;
        RECT 91.860 177.700 94.060 179.110 ;
        RECT 95.220 177.700 97.420 179.110 ;
        RECT 98.580 177.700 100.780 179.110 ;
        RECT 101.940 177.700 104.140 179.110 ;
        RECT 105.300 177.700 108.620 179.110 ;
        RECT 109.780 177.700 111.980 179.110 ;
        RECT 113.140 177.700 115.340 179.110 ;
        RECT 116.500 177.700 118.700 179.110 ;
        RECT 119.860 177.700 122.060 179.110 ;
        RECT 123.220 177.700 126.540 179.110 ;
        RECT 127.700 177.700 129.900 179.110 ;
        RECT 131.060 177.700 133.260 179.110 ;
        RECT 134.420 177.700 136.620 179.110 ;
        RECT 137.780 177.700 139.980 179.110 ;
        RECT 141.140 177.700 144.460 179.110 ;
        RECT 145.620 177.700 147.820 179.110 ;
        RECT 148.980 177.700 151.180 179.110 ;
        RECT 152.340 177.700 154.540 179.110 ;
        RECT 155.700 177.700 157.900 179.110 ;
        RECT 159.060 177.700 162.380 179.110 ;
        RECT 163.540 177.700 165.740 179.110 ;
        RECT 166.900 177.700 169.100 179.110 ;
        RECT 170.260 177.700 172.460 179.110 ;
        RECT 173.620 177.700 175.820 179.110 ;
        RECT 176.980 177.700 180.300 179.110 ;
        RECT 181.460 177.700 183.660 179.110 ;
        RECT 184.820 177.700 187.020 179.110 ;
        RECT 188.180 177.700 190.380 179.110 ;
        RECT 191.540 177.700 193.740 179.110 ;
        RECT 194.900 177.700 198.220 179.110 ;
        RECT 199.380 177.700 201.580 179.110 ;
        RECT 202.740 177.700 204.940 179.110 ;
        RECT 206.100 177.700 208.300 179.110 ;
        RECT 209.460 177.700 211.660 179.110 ;
        RECT 212.820 177.700 216.140 179.110 ;
        RECT 217.300 177.700 219.500 179.110 ;
        RECT 220.660 177.700 222.860 179.110 ;
        RECT 224.020 177.700 226.220 179.110 ;
        RECT 227.380 177.700 229.580 179.110 ;
        RECT 230.740 177.700 234.060 179.110 ;
        RECT 235.220 177.700 237.420 179.110 ;
        RECT 238.580 177.700 240.780 179.110 ;
        RECT 241.940 177.700 244.140 179.110 ;
        RECT 245.300 177.700 247.500 179.110 ;
        RECT 248.660 177.700 251.980 179.110 ;
        RECT 253.140 177.700 255.340 179.110 ;
        RECT 256.500 177.700 258.700 179.110 ;
        RECT 259.860 177.700 262.060 179.110 ;
        RECT 263.220 177.700 265.420 179.110 ;
        RECT 266.580 177.700 269.900 179.110 ;
        RECT 271.060 177.700 273.260 179.110 ;
        RECT 274.420 177.700 276.620 179.110 ;
        RECT 277.780 177.700 279.980 179.110 ;
        RECT 281.140 177.700 283.340 179.110 ;
        RECT 284.500 177.700 287.820 179.110 ;
        RECT 288.980 177.700 291.180 179.110 ;
        RECT 292.340 177.700 294.540 179.110 ;
        RECT 295.700 177.700 297.900 179.110 ;
        RECT 299.060 177.700 301.260 179.110 ;
        RECT 302.420 177.700 305.740 179.110 ;
        RECT 306.900 177.700 309.100 179.110 ;
        RECT 310.260 177.700 312.460 179.110 ;
        RECT 313.620 177.700 315.820 179.110 ;
        RECT 316.980 177.700 319.180 179.110 ;
        RECT 320.340 177.700 323.660 179.110 ;
        RECT 324.820 177.700 327.020 179.110 ;
        RECT 328.180 177.700 330.380 179.110 ;
        RECT 331.540 177.700 333.740 179.110 ;
        RECT 334.900 177.700 337.100 179.110 ;
        RECT 338.260 177.700 341.580 179.110 ;
        RECT 342.740 177.700 344.940 179.110 ;
        RECT 346.100 177.700 348.300 179.110 ;
        RECT 349.460 177.700 351.660 179.110 ;
        RECT 352.820 177.700 355.020 179.110 ;
        RECT 356.180 177.700 359.500 179.110 ;
        RECT 360.660 177.700 362.860 179.110 ;
        RECT 364.020 177.700 366.220 179.110 ;
        RECT 367.380 177.700 369.580 179.110 ;
        RECT 370.740 177.700 372.940 179.110 ;
        RECT 374.100 177.700 377.420 179.110 ;
        RECT 378.580 177.700 380.780 179.110 ;
        RECT 381.940 177.700 384.140 179.110 ;
        RECT 385.300 177.700 387.500 179.110 ;
        RECT 388.660 177.700 390.860 179.110 ;
        RECT 392.020 177.700 395.340 179.110 ;
        RECT 396.500 177.700 398.700 179.110 ;
        RECT 399.860 177.700 402.060 179.110 ;
        RECT 403.220 177.700 405.420 179.110 ;
        RECT 406.580 177.700 408.780 179.110 ;
        RECT 409.940 177.700 413.260 179.110 ;
        RECT 414.420 177.700 416.620 179.110 ;
        RECT 417.780 177.700 419.980 179.110 ;
        RECT 421.140 177.700 423.340 179.110 ;
        RECT 424.500 177.700 426.700 179.110 ;
        RECT 427.860 177.700 431.180 179.110 ;
        RECT 432.340 177.700 434.540 179.110 ;
        RECT 435.700 177.700 437.900 179.110 ;
        RECT 439.060 177.700 441.260 179.110 ;
        RECT 442.420 177.700 444.620 179.110 ;
        RECT 1.820 2.300 445.060 177.700 ;
        RECT 2.260 1.400 22.380 2.300 ;
        RECT 23.540 1.400 43.660 2.300 ;
        RECT 44.820 1.400 64.940 2.300 ;
        RECT 66.100 1.400 86.220 2.300 ;
        RECT 87.380 1.400 107.500 2.300 ;
        RECT 108.660 1.400 128.780 2.300 ;
        RECT 129.940 1.400 150.060 2.300 ;
        RECT 151.220 1.400 171.340 2.300 ;
        RECT 172.500 1.400 192.620 2.300 ;
        RECT 193.780 1.400 213.900 2.300 ;
        RECT 215.060 1.400 235.180 2.300 ;
        RECT 236.340 1.400 256.460 2.300 ;
        RECT 257.620 1.400 277.740 2.300 ;
        RECT 278.900 1.400 299.020 2.300 ;
        RECT 300.180 1.400 320.300 2.300 ;
        RECT 321.460 1.400 341.580 2.300 ;
        RECT 342.740 1.400 362.860 2.300 ;
        RECT 364.020 1.400 384.140 2.300 ;
        RECT 385.300 1.400 405.420 2.300 ;
        RECT 406.580 1.400 426.700 2.300 ;
        RECT 427.860 1.400 445.060 2.300 ;
      LAYER Metal3 ;
        RECT 1.770 7.700 445.110 179.060 ;
  END
END S_term_single2
END LIBRARY

