VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO N_term_single
  CLASS BLOCK ;
  FOREIGN N_term_single ;
  ORIGIN 0.000 0.000 ;
  SIZE 390.000 BY 180.000 ;
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.560 0.000 162.120 2.000 ;
    END
  END Ci
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 327.320 0.000 327.880 2.000 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 358.680 0.000 359.240 2.000 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 362.040 0.000 362.600 2.000 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 364.280 0.000 364.840 2.000 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 367.640 0.000 368.200 2.000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 371.000 0.000 371.560 2.000 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 374.360 0.000 374.920 2.000 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 376.600 0.000 377.160 2.000 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 379.960 0.000 380.520 2.000 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 383.320 0.000 383.880 2.000 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.680 0.000 387.240 2.000 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 330.680 0.000 331.240 2.000 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 334.040 0.000 334.600 2.000 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 337.400 0.000 337.960 2.000 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 339.640 0.000 340.200 2.000 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 343.000 0.000 343.560 2.000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 346.360 0.000 346.920 2.000 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 349.720 0.000 350.280 2.000 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 351.960 0.000 352.520 2.000 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 355.320 0.000 355.880 2.000 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 19.320 178.000 19.880 180.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.120 178.000 204.680 180.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 223.160 178.000 223.720 180.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.080 178.000 241.640 180.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 260.120 178.000 260.680 180.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.040 178.000 278.600 180.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 297.080 178.000 297.640 180.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.000 178.000 315.560 180.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 334.040 178.000 334.600 180.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 351.960 178.000 352.520 180.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 371.000 178.000 371.560 180.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 38.360 178.000 38.920 180.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 56.280 178.000 56.840 180.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 75.320 178.000 75.880 180.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 93.240 178.000 93.800 180.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 112.280 178.000 112.840 180.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 130.200 178.000 130.760 180.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 149.240 178.000 149.800 180.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 167.160 178.000 167.720 180.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 186.200 178.000 186.760 180.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1.400 0.000 1.960 2.000 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.640 0.000 4.200 2.000 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 7.000 0.000 7.560 2.000 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.360 0.000 10.920 2.000 ;
    END
  END N1END[3]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 38.360 0.000 38.920 2.000 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.600 0.000 41.160 2.000 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.960 0.000 44.520 2.000 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.320 0.000 47.880 2.000 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.680 0.000 51.240 2.000 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 52.920 0.000 53.480 2.000 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 56.280 0.000 56.840 2.000 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 59.640 0.000 60.200 2.000 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.720 0.000 14.280 2.000 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 15.960 0.000 16.520 2.000 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 19.320 0.000 19.880 2.000 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 22.680 0.000 23.240 2.000 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.040 0.000 26.600 2.000 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 28.280 0.000 28.840 2.000 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 31.640 0.000 32.200 2.000 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 35.000 0.000 35.560 2.000 ;
    END
  END N2MID[7]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.000 0.000 63.560 2.000 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 93.240 0.000 93.800 2.000 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 96.600 0.000 97.160 2.000 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 99.960 0.000 100.520 2.000 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 102.200 0.000 102.760 2.000 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 105.560 0.000 106.120 2.000 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 108.920 0.000 109.480 2.000 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 65.240 0.000 65.800 2.000 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 68.600 0.000 69.160 2.000 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 71.960 0.000 72.520 2.000 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 75.320 0.000 75.880 2.000 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.560 0.000 78.120 2.000 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.920 0.000 81.480 2.000 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.280 0.000 84.840 2.000 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.640 0.000 88.200 2.000 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 89.880 0.000 90.440 2.000 ;
    END
  END N4END[9]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 112.280 0.000 112.840 2.000 ;
    END
  END NN4END[0]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 142.520 0.000 143.080 2.000 ;
    END
  END NN4END[10]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 145.880 0.000 146.440 2.000 ;
    END
  END NN4END[11]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 149.240 0.000 149.800 2.000 ;
    END
  END NN4END[12]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.480 0.000 152.040 2.000 ;
    END
  END NN4END[13]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.840 0.000 155.400 2.000 ;
    END
  END NN4END[14]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 158.200 0.000 158.760 2.000 ;
    END
  END NN4END[15]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 114.520 0.000 115.080 2.000 ;
    END
  END NN4END[1]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.880 0.000 118.440 2.000 ;
    END
  END NN4END[2]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 121.240 0.000 121.800 2.000 ;
    END
  END NN4END[3]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.600 0.000 125.160 2.000 ;
    END
  END NN4END[4]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 126.840 0.000 127.400 2.000 ;
    END
  END NN4END[5]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 130.200 0.000 130.760 2.000 ;
    END
  END NN4END[6]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 133.560 0.000 134.120 2.000 ;
    END
  END NN4END[7]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 136.920 0.000 137.480 2.000 ;
    END
  END NN4END[8]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 139.160 0.000 139.720 2.000 ;
    END
  END NN4END[9]
  PIN S1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 163.800 0.000 164.360 2.000 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 167.160 0.000 167.720 2.000 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 170.520 0.000 171.080 2.000 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 173.880 0.000 174.440 2.000 ;
    END
  END S1BEG[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 176.120 0.000 176.680 2.000 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 179.480 0.000 180.040 2.000 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 182.840 0.000 183.400 2.000 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 186.200 0.000 186.760 2.000 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 188.440 0.000 189.000 2.000 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 191.800 0.000 192.360 2.000 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 195.160 0.000 195.720 2.000 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 198.520 0.000 199.080 2.000 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.880 0.000 202.440 2.000 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.120 0.000 204.680 2.000 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 207.480 0.000 208.040 2.000 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 210.840 0.000 211.400 2.000 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 214.200 0.000 214.760 2.000 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 216.440 0.000 217.000 2.000 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 219.800 0.000 220.360 2.000 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 223.160 0.000 223.720 2.000 ;
    END
  END S2BEGb[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 226.520 0.000 227.080 2.000 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 256.760 0.000 257.320 2.000 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 260.120 0.000 260.680 2.000 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 263.480 0.000 264.040 2.000 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 265.720 0.000 266.280 2.000 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 269.080 0.000 269.640 2.000 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 272.440 0.000 273.000 2.000 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.760 0.000 229.320 2.000 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 232.120 0.000 232.680 2.000 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 235.480 0.000 236.040 2.000 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.840 0.000 239.400 2.000 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.080 0.000 241.640 2.000 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 244.440 0.000 245.000 2.000 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 247.800 0.000 248.360 2.000 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 251.160 0.000 251.720 2.000 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 253.400 0.000 253.960 2.000 ;
    END
  END S4BEG[9]
  PIN SS4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.800 0.000 276.360 2.000 ;
    END
  END SS4BEG[0]
  PIN SS4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 306.040 0.000 306.600 2.000 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 309.400 0.000 309.960 2.000 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 312.760 0.000 313.320 2.000 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.000 0.000 315.560 2.000 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 318.360 0.000 318.920 2.000 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 321.720 0.000 322.280 2.000 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.040 0.000 278.600 2.000 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 281.400 0.000 281.960 2.000 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 284.760 0.000 285.320 2.000 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.120 0.000 288.680 2.000 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 290.360 0.000 290.920 2.000 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 293.720 0.000 294.280 2.000 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 297.080 0.000 297.640 2.000 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 300.440 0.000 301.000 2.000 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.680 0.000 303.240 2.000 ;
    END
  END SS4BEG[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 325.080 0.000 325.640 2.000 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1.400 178.000 1.960 180.000 ;
    END
  END UserCLKo
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 52.960 7.540 54.560 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 147.040 7.540 148.640 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 241.120 7.540 242.720 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 335.200 7.540 336.800 168.860 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 100.000 7.540 101.600 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 194.080 7.540 195.680 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 288.160 7.540 289.760 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 382.240 7.540 383.840 168.860 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 6.720 6.870 383.840 168.860 ;
      LAYER Metal2 ;
        RECT 2.260 177.700 19.020 178.500 ;
        RECT 20.180 177.700 38.060 178.500 ;
        RECT 39.220 177.700 55.980 178.500 ;
        RECT 57.140 177.700 75.020 178.500 ;
        RECT 76.180 177.700 92.940 178.500 ;
        RECT 94.100 177.700 111.980 178.500 ;
        RECT 113.140 177.700 129.900 178.500 ;
        RECT 131.060 177.700 148.940 178.500 ;
        RECT 150.100 177.700 166.860 178.500 ;
        RECT 168.020 177.700 185.900 178.500 ;
        RECT 187.060 177.700 203.820 178.500 ;
        RECT 204.980 177.700 222.860 178.500 ;
        RECT 224.020 177.700 240.780 178.500 ;
        RECT 241.940 177.700 259.820 178.500 ;
        RECT 260.980 177.700 277.740 178.500 ;
        RECT 278.900 177.700 296.780 178.500 ;
        RECT 297.940 177.700 314.700 178.500 ;
        RECT 315.860 177.700 333.740 178.500 ;
        RECT 334.900 177.700 351.660 178.500 ;
        RECT 352.820 177.700 370.700 178.500 ;
        RECT 371.860 177.700 386.820 178.500 ;
        RECT 1.820 2.300 386.820 177.700 ;
        RECT 2.260 1.260 3.340 2.300 ;
        RECT 4.500 1.260 6.700 2.300 ;
        RECT 7.860 1.260 10.060 2.300 ;
        RECT 11.220 1.260 13.420 2.300 ;
        RECT 14.580 1.260 15.660 2.300 ;
        RECT 16.820 1.260 19.020 2.300 ;
        RECT 20.180 1.260 22.380 2.300 ;
        RECT 23.540 1.260 25.740 2.300 ;
        RECT 26.900 1.260 27.980 2.300 ;
        RECT 29.140 1.260 31.340 2.300 ;
        RECT 32.500 1.260 34.700 2.300 ;
        RECT 35.860 1.260 38.060 2.300 ;
        RECT 39.220 1.260 40.300 2.300 ;
        RECT 41.460 1.260 43.660 2.300 ;
        RECT 44.820 1.260 47.020 2.300 ;
        RECT 48.180 1.260 50.380 2.300 ;
        RECT 51.540 1.260 52.620 2.300 ;
        RECT 53.780 1.260 55.980 2.300 ;
        RECT 57.140 1.260 59.340 2.300 ;
        RECT 60.500 1.260 62.700 2.300 ;
        RECT 63.860 1.260 64.940 2.300 ;
        RECT 66.100 1.260 68.300 2.300 ;
        RECT 69.460 1.260 71.660 2.300 ;
        RECT 72.820 1.260 75.020 2.300 ;
        RECT 76.180 1.260 77.260 2.300 ;
        RECT 78.420 1.260 80.620 2.300 ;
        RECT 81.780 1.260 83.980 2.300 ;
        RECT 85.140 1.260 87.340 2.300 ;
        RECT 88.500 1.260 89.580 2.300 ;
        RECT 90.740 1.260 92.940 2.300 ;
        RECT 94.100 1.260 96.300 2.300 ;
        RECT 97.460 1.260 99.660 2.300 ;
        RECT 100.820 1.260 101.900 2.300 ;
        RECT 103.060 1.260 105.260 2.300 ;
        RECT 106.420 1.260 108.620 2.300 ;
        RECT 109.780 1.260 111.980 2.300 ;
        RECT 113.140 1.260 114.220 2.300 ;
        RECT 115.380 1.260 117.580 2.300 ;
        RECT 118.740 1.260 120.940 2.300 ;
        RECT 122.100 1.260 124.300 2.300 ;
        RECT 125.460 1.260 126.540 2.300 ;
        RECT 127.700 1.260 129.900 2.300 ;
        RECT 131.060 1.260 133.260 2.300 ;
        RECT 134.420 1.260 136.620 2.300 ;
        RECT 137.780 1.260 138.860 2.300 ;
        RECT 140.020 1.260 142.220 2.300 ;
        RECT 143.380 1.260 145.580 2.300 ;
        RECT 146.740 1.260 148.940 2.300 ;
        RECT 150.100 1.260 151.180 2.300 ;
        RECT 152.340 1.260 154.540 2.300 ;
        RECT 155.700 1.260 157.900 2.300 ;
        RECT 159.060 1.260 161.260 2.300 ;
        RECT 162.420 1.260 163.500 2.300 ;
        RECT 164.660 1.260 166.860 2.300 ;
        RECT 168.020 1.260 170.220 2.300 ;
        RECT 171.380 1.260 173.580 2.300 ;
        RECT 174.740 1.260 175.820 2.300 ;
        RECT 176.980 1.260 179.180 2.300 ;
        RECT 180.340 1.260 182.540 2.300 ;
        RECT 183.700 1.260 185.900 2.300 ;
        RECT 187.060 1.260 188.140 2.300 ;
        RECT 189.300 1.260 191.500 2.300 ;
        RECT 192.660 1.260 194.860 2.300 ;
        RECT 196.020 1.260 198.220 2.300 ;
        RECT 199.380 1.260 201.580 2.300 ;
        RECT 202.740 1.260 203.820 2.300 ;
        RECT 204.980 1.260 207.180 2.300 ;
        RECT 208.340 1.260 210.540 2.300 ;
        RECT 211.700 1.260 213.900 2.300 ;
        RECT 215.060 1.260 216.140 2.300 ;
        RECT 217.300 1.260 219.500 2.300 ;
        RECT 220.660 1.260 222.860 2.300 ;
        RECT 224.020 1.260 226.220 2.300 ;
        RECT 227.380 1.260 228.460 2.300 ;
        RECT 229.620 1.260 231.820 2.300 ;
        RECT 232.980 1.260 235.180 2.300 ;
        RECT 236.340 1.260 238.540 2.300 ;
        RECT 239.700 1.260 240.780 2.300 ;
        RECT 241.940 1.260 244.140 2.300 ;
        RECT 245.300 1.260 247.500 2.300 ;
        RECT 248.660 1.260 250.860 2.300 ;
        RECT 252.020 1.260 253.100 2.300 ;
        RECT 254.260 1.260 256.460 2.300 ;
        RECT 257.620 1.260 259.820 2.300 ;
        RECT 260.980 1.260 263.180 2.300 ;
        RECT 264.340 1.260 265.420 2.300 ;
        RECT 266.580 1.260 268.780 2.300 ;
        RECT 269.940 1.260 272.140 2.300 ;
        RECT 273.300 1.260 275.500 2.300 ;
        RECT 276.660 1.260 277.740 2.300 ;
        RECT 278.900 1.260 281.100 2.300 ;
        RECT 282.260 1.260 284.460 2.300 ;
        RECT 285.620 1.260 287.820 2.300 ;
        RECT 288.980 1.260 290.060 2.300 ;
        RECT 291.220 1.260 293.420 2.300 ;
        RECT 294.580 1.260 296.780 2.300 ;
        RECT 297.940 1.260 300.140 2.300 ;
        RECT 301.300 1.260 302.380 2.300 ;
        RECT 303.540 1.260 305.740 2.300 ;
        RECT 306.900 1.260 309.100 2.300 ;
        RECT 310.260 1.260 312.460 2.300 ;
        RECT 313.620 1.260 314.700 2.300 ;
        RECT 315.860 1.260 318.060 2.300 ;
        RECT 319.220 1.260 321.420 2.300 ;
        RECT 322.580 1.260 324.780 2.300 ;
        RECT 325.940 1.260 327.020 2.300 ;
        RECT 328.180 1.260 330.380 2.300 ;
        RECT 331.540 1.260 333.740 2.300 ;
        RECT 334.900 1.260 337.100 2.300 ;
        RECT 338.260 1.260 339.340 2.300 ;
        RECT 340.500 1.260 342.700 2.300 ;
        RECT 343.860 1.260 346.060 2.300 ;
        RECT 347.220 1.260 349.420 2.300 ;
        RECT 350.580 1.260 351.660 2.300 ;
        RECT 352.820 1.260 355.020 2.300 ;
        RECT 356.180 1.260 358.380 2.300 ;
        RECT 359.540 1.260 361.740 2.300 ;
        RECT 362.900 1.260 363.980 2.300 ;
        RECT 365.140 1.260 367.340 2.300 ;
        RECT 368.500 1.260 370.700 2.300 ;
        RECT 371.860 1.260 374.060 2.300 ;
        RECT 375.220 1.260 376.300 2.300 ;
        RECT 377.460 1.260 379.660 2.300 ;
        RECT 380.820 1.260 383.020 2.300 ;
        RECT 384.180 1.260 386.380 2.300 ;
      LAYER Metal3 ;
        RECT 1.770 2.940 386.870 168.700 ;
      LAYER Metal4 ;
        RECT 141.260 12.970 146.740 30.710 ;
        RECT 148.940 12.970 193.780 30.710 ;
        RECT 195.980 12.970 234.500 30.710 ;
  END
END N_term_single
END LIBRARY

