VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO N_term_single2
  CLASS BLOCK ;
  FOREIGN N_term_single2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 450.000 BY 180.000 ;
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 377.720 0.000 378.280 2.000 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 413.560 0.000 414.120 2.000 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 416.920 0.000 417.480 2.000 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 420.280 0.000 420.840 2.000 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 423.640 0.000 424.200 2.000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 427.000 0.000 427.560 2.000 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 431.480 0.000 432.040 2.000 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 434.840 0.000 435.400 2.000 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 438.200 0.000 438.760 2.000 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 441.560 0.000 442.120 2.000 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 444.920 0.000 445.480 2.000 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 381.080 0.000 381.640 2.000 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 384.440 0.000 385.000 2.000 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 387.800 0.000 388.360 2.000 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 391.160 0.000 391.720 2.000 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 395.640 0.000 396.200 2.000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 399.000 0.000 399.560 2.000 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 402.360 0.000 402.920 2.000 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 405.720 0.000 406.280 2.000 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 409.080 0.000 409.640 2.000 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 22.680 178.000 23.240 180.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 235.480 178.000 236.040 180.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 256.760 178.000 257.320 180.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.040 178.000 278.600 180.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 299.320 178.000 299.880 180.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 320.600 178.000 321.160 180.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 341.880 178.000 342.440 180.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 363.160 178.000 363.720 180.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 384.440 178.000 385.000 180.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 405.720 178.000 406.280 180.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 427.000 178.000 427.560 180.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.960 178.000 44.520 180.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 65.240 178.000 65.800 180.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 86.520 178.000 87.080 180.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.800 178.000 108.360 180.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 129.080 178.000 129.640 180.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 150.360 178.000 150.920 180.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.640 178.000 172.200 180.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 192.920 178.000 193.480 180.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 214.200 178.000 214.760 180.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1.400 0.000 1.960 2.000 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 4.760 0.000 5.320 2.000 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 8.120 0.000 8.680 2.000 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 11.480 0.000 12.040 2.000 ;
    END
  END N1END[3]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.960 0.000 44.520 2.000 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.320 0.000 47.880 2.000 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.680 0.000 51.240 2.000 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 55.160 0.000 55.720 2.000 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 58.520 0.000 59.080 2.000 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 61.880 0.000 62.440 2.000 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 65.240 0.000 65.800 2.000 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 68.600 0.000 69.160 2.000 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 14.840 0.000 15.400 2.000 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 19.320 0.000 19.880 2.000 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 22.680 0.000 23.240 2.000 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.040 0.000 26.600 2.000 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 29.400 0.000 29.960 2.000 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 32.760 0.000 33.320 2.000 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 37.240 0.000 37.800 2.000 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.600 0.000 41.160 2.000 ;
    END
  END N2MID[7]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.080 0.000 73.640 2.000 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 108.920 0.000 109.480 2.000 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 112.280 0.000 112.840 2.000 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 115.640 0.000 116.200 2.000 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 119.000 0.000 119.560 2.000 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 122.360 0.000 122.920 2.000 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 126.840 0.000 127.400 2.000 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 76.440 0.000 77.000 2.000 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 79.800 0.000 80.360 2.000 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 83.160 0.000 83.720 2.000 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 86.520 0.000 87.080 2.000 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 91.000 0.000 91.560 2.000 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.360 0.000 94.920 2.000 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.720 0.000 98.280 2.000 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 101.080 0.000 101.640 2.000 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.440 0.000 105.000 2.000 ;
    END
  END N4END[9]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 130.200 0.000 130.760 2.000 ;
    END
  END NN4END[0]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 166.040 0.000 166.600 2.000 ;
    END
  END NN4END[10]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 169.400 0.000 169.960 2.000 ;
    END
  END NN4END[11]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 172.760 0.000 173.320 2.000 ;
    END
  END NN4END[12]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 176.120 0.000 176.680 2.000 ;
    END
  END NN4END[13]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 180.600 0.000 181.160 2.000 ;
    END
  END NN4END[14]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 183.960 0.000 184.520 2.000 ;
    END
  END NN4END[15]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 133.560 0.000 134.120 2.000 ;
    END
  END NN4END[1]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 136.920 0.000 137.480 2.000 ;
    END
  END NN4END[2]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 140.280 0.000 140.840 2.000 ;
    END
  END NN4END[3]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.760 0.000 145.320 2.000 ;
    END
  END NN4END[4]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 148.120 0.000 148.680 2.000 ;
    END
  END NN4END[5]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.480 0.000 152.040 2.000 ;
    END
  END NN4END[6]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.840 0.000 155.400 2.000 ;
    END
  END NN4END[7]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 158.200 0.000 158.760 2.000 ;
    END
  END NN4END[8]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 162.680 0.000 163.240 2.000 ;
    END
  END NN4END[9]
  PIN S1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 187.320 0.000 187.880 2.000 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 190.680 0.000 191.240 2.000 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.040 0.000 194.600 2.000 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 198.520 0.000 199.080 2.000 ;
    END
  END S1BEG[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.880 0.000 202.440 2.000 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 205.240 0.000 205.800 2.000 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 208.600 0.000 209.160 2.000 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.960 0.000 212.520 2.000 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 216.440 0.000 217.000 2.000 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 219.800 0.000 220.360 2.000 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 223.160 0.000 223.720 2.000 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 226.520 0.000 227.080 2.000 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 229.880 0.000 230.440 2.000 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.360 0.000 234.920 2.000 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 237.720 0.000 238.280 2.000 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.080 0.000 241.640 2.000 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 244.440 0.000 245.000 2.000 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 247.800 0.000 248.360 2.000 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 252.280 0.000 252.840 2.000 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 255.640 0.000 256.200 2.000 ;
    END
  END S2BEGb[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 259.000 0.000 259.560 2.000 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 294.840 0.000 295.400 2.000 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 298.200 0.000 298.760 2.000 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 301.560 0.000 302.120 2.000 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 306.040 0.000 306.600 2.000 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 309.400 0.000 309.960 2.000 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 312.760 0.000 313.320 2.000 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.360 0.000 262.920 2.000 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 265.720 0.000 266.280 2.000 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 270.200 0.000 270.760 2.000 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 273.560 0.000 274.120 2.000 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 276.920 0.000 277.480 2.000 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 280.280 0.000 280.840 2.000 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 283.640 0.000 284.200 2.000 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.120 0.000 288.680 2.000 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 291.480 0.000 292.040 2.000 ;
    END
  END S4BEG[9]
  PIN SS4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 316.120 0.000 316.680 2.000 ;
    END
  END SS4BEG[0]
  PIN SS4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 351.960 0.000 352.520 2.000 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 355.320 0.000 355.880 2.000 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 359.800 0.000 360.360 2.000 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 363.160 0.000 363.720 2.000 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 366.520 0.000 367.080 2.000 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 369.880 0.000 370.440 2.000 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 319.480 0.000 320.040 2.000 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 323.960 0.000 324.520 2.000 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 327.320 0.000 327.880 2.000 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 330.680 0.000 331.240 2.000 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 334.040 0.000 334.600 2.000 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 337.400 0.000 337.960 2.000 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 341.880 0.000 342.440 2.000 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 345.240 0.000 345.800 2.000 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 348.600 0.000 349.160 2.000 ;
    END
  END SS4BEG[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 373.240 0.000 373.800 2.000 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1.400 178.000 1.960 180.000 ;
    END
  END UserCLKo
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 60.445 7.540 62.045 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 169.500 7.540 171.100 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 278.555 7.540 280.155 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 387.610 7.540 389.210 168.860 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 114.970 7.540 116.570 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 224.025 7.540 225.625 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 333.080 7.540 334.680 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 442.135 7.540 443.735 168.860 ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        RECT 6.720 7.540 443.735 168.860 ;
      LAYER Metal2 ;
        RECT 2.260 177.700 22.380 178.500 ;
        RECT 23.540 177.700 43.660 178.500 ;
        RECT 44.820 177.700 64.940 178.500 ;
        RECT 66.100 177.700 86.220 178.500 ;
        RECT 87.380 177.700 107.500 178.500 ;
        RECT 108.660 177.700 128.780 178.500 ;
        RECT 129.940 177.700 150.060 178.500 ;
        RECT 151.220 177.700 171.340 178.500 ;
        RECT 172.500 177.700 192.620 178.500 ;
        RECT 193.780 177.700 213.900 178.500 ;
        RECT 215.060 177.700 235.180 178.500 ;
        RECT 236.340 177.700 256.460 178.500 ;
        RECT 257.620 177.700 277.740 178.500 ;
        RECT 278.900 177.700 299.020 178.500 ;
        RECT 300.180 177.700 320.300 178.500 ;
        RECT 321.460 177.700 341.580 178.500 ;
        RECT 342.740 177.700 362.860 178.500 ;
        RECT 364.020 177.700 384.140 178.500 ;
        RECT 385.300 177.700 405.420 178.500 ;
        RECT 406.580 177.700 426.700 178.500 ;
        RECT 427.860 177.700 445.060 178.500 ;
        RECT 1.820 2.300 445.060 177.700 ;
        RECT 2.260 1.260 4.460 2.300 ;
        RECT 5.620 1.260 7.820 2.300 ;
        RECT 8.980 1.260 11.180 2.300 ;
        RECT 12.340 1.260 14.540 2.300 ;
        RECT 15.700 1.260 19.020 2.300 ;
        RECT 20.180 1.260 22.380 2.300 ;
        RECT 23.540 1.260 25.740 2.300 ;
        RECT 26.900 1.260 29.100 2.300 ;
        RECT 30.260 1.260 32.460 2.300 ;
        RECT 33.620 1.260 36.940 2.300 ;
        RECT 38.100 1.260 40.300 2.300 ;
        RECT 41.460 1.260 43.660 2.300 ;
        RECT 44.820 1.260 47.020 2.300 ;
        RECT 48.180 1.260 50.380 2.300 ;
        RECT 51.540 1.260 54.860 2.300 ;
        RECT 56.020 1.260 58.220 2.300 ;
        RECT 59.380 1.260 61.580 2.300 ;
        RECT 62.740 1.260 64.940 2.300 ;
        RECT 66.100 1.260 68.300 2.300 ;
        RECT 69.460 1.260 72.780 2.300 ;
        RECT 73.940 1.260 76.140 2.300 ;
        RECT 77.300 1.260 79.500 2.300 ;
        RECT 80.660 1.260 82.860 2.300 ;
        RECT 84.020 1.260 86.220 2.300 ;
        RECT 87.380 1.260 90.700 2.300 ;
        RECT 91.860 1.260 94.060 2.300 ;
        RECT 95.220 1.260 97.420 2.300 ;
        RECT 98.580 1.260 100.780 2.300 ;
        RECT 101.940 1.260 104.140 2.300 ;
        RECT 105.300 1.260 108.620 2.300 ;
        RECT 109.780 1.260 111.980 2.300 ;
        RECT 113.140 1.260 115.340 2.300 ;
        RECT 116.500 1.260 118.700 2.300 ;
        RECT 119.860 1.260 122.060 2.300 ;
        RECT 123.220 1.260 126.540 2.300 ;
        RECT 127.700 1.260 129.900 2.300 ;
        RECT 131.060 1.260 133.260 2.300 ;
        RECT 134.420 1.260 136.620 2.300 ;
        RECT 137.780 1.260 139.980 2.300 ;
        RECT 141.140 1.260 144.460 2.300 ;
        RECT 145.620 1.260 147.820 2.300 ;
        RECT 148.980 1.260 151.180 2.300 ;
        RECT 152.340 1.260 154.540 2.300 ;
        RECT 155.700 1.260 157.900 2.300 ;
        RECT 159.060 1.260 162.380 2.300 ;
        RECT 163.540 1.260 165.740 2.300 ;
        RECT 166.900 1.260 169.100 2.300 ;
        RECT 170.260 1.260 172.460 2.300 ;
        RECT 173.620 1.260 175.820 2.300 ;
        RECT 176.980 1.260 180.300 2.300 ;
        RECT 181.460 1.260 183.660 2.300 ;
        RECT 184.820 1.260 187.020 2.300 ;
        RECT 188.180 1.260 190.380 2.300 ;
        RECT 191.540 1.260 193.740 2.300 ;
        RECT 194.900 1.260 198.220 2.300 ;
        RECT 199.380 1.260 201.580 2.300 ;
        RECT 202.740 1.260 204.940 2.300 ;
        RECT 206.100 1.260 208.300 2.300 ;
        RECT 209.460 1.260 211.660 2.300 ;
        RECT 212.820 1.260 216.140 2.300 ;
        RECT 217.300 1.260 219.500 2.300 ;
        RECT 220.660 1.260 222.860 2.300 ;
        RECT 224.020 1.260 226.220 2.300 ;
        RECT 227.380 1.260 229.580 2.300 ;
        RECT 230.740 1.260 234.060 2.300 ;
        RECT 235.220 1.260 237.420 2.300 ;
        RECT 238.580 1.260 240.780 2.300 ;
        RECT 241.940 1.260 244.140 2.300 ;
        RECT 245.300 1.260 247.500 2.300 ;
        RECT 248.660 1.260 251.980 2.300 ;
        RECT 253.140 1.260 255.340 2.300 ;
        RECT 256.500 1.260 258.700 2.300 ;
        RECT 259.860 1.260 262.060 2.300 ;
        RECT 263.220 1.260 265.420 2.300 ;
        RECT 266.580 1.260 269.900 2.300 ;
        RECT 271.060 1.260 273.260 2.300 ;
        RECT 274.420 1.260 276.620 2.300 ;
        RECT 277.780 1.260 279.980 2.300 ;
        RECT 281.140 1.260 283.340 2.300 ;
        RECT 284.500 1.260 287.820 2.300 ;
        RECT 288.980 1.260 291.180 2.300 ;
        RECT 292.340 1.260 294.540 2.300 ;
        RECT 295.700 1.260 297.900 2.300 ;
        RECT 299.060 1.260 301.260 2.300 ;
        RECT 302.420 1.260 305.740 2.300 ;
        RECT 306.900 1.260 309.100 2.300 ;
        RECT 310.260 1.260 312.460 2.300 ;
        RECT 313.620 1.260 315.820 2.300 ;
        RECT 316.980 1.260 319.180 2.300 ;
        RECT 320.340 1.260 323.660 2.300 ;
        RECT 324.820 1.260 327.020 2.300 ;
        RECT 328.180 1.260 330.380 2.300 ;
        RECT 331.540 1.260 333.740 2.300 ;
        RECT 334.900 1.260 337.100 2.300 ;
        RECT 338.260 1.260 341.580 2.300 ;
        RECT 342.740 1.260 344.940 2.300 ;
        RECT 346.100 1.260 348.300 2.300 ;
        RECT 349.460 1.260 351.660 2.300 ;
        RECT 352.820 1.260 355.020 2.300 ;
        RECT 356.180 1.260 359.500 2.300 ;
        RECT 360.660 1.260 362.860 2.300 ;
        RECT 364.020 1.260 366.220 2.300 ;
        RECT 367.380 1.260 369.580 2.300 ;
        RECT 370.740 1.260 372.940 2.300 ;
        RECT 374.100 1.260 377.420 2.300 ;
        RECT 378.580 1.260 380.780 2.300 ;
        RECT 381.940 1.260 384.140 2.300 ;
        RECT 385.300 1.260 387.500 2.300 ;
        RECT 388.660 1.260 390.860 2.300 ;
        RECT 392.020 1.260 395.340 2.300 ;
        RECT 396.500 1.260 398.700 2.300 ;
        RECT 399.860 1.260 402.060 2.300 ;
        RECT 403.220 1.260 405.420 2.300 ;
        RECT 406.580 1.260 408.780 2.300 ;
        RECT 409.940 1.260 413.260 2.300 ;
        RECT 414.420 1.260 416.620 2.300 ;
        RECT 417.780 1.260 419.980 2.300 ;
        RECT 421.140 1.260 423.340 2.300 ;
        RECT 424.500 1.260 426.700 2.300 ;
        RECT 427.860 1.260 431.180 2.300 ;
        RECT 432.340 1.260 434.540 2.300 ;
        RECT 435.700 1.260 437.900 2.300 ;
        RECT 439.060 1.260 441.260 2.300 ;
        RECT 442.420 1.260 444.620 2.300 ;
      LAYER Metal3 ;
        RECT 1.770 2.380 445.110 168.700 ;
      LAYER Metal4 ;
        RECT 129.500 8.490 169.200 27.910 ;
        RECT 171.400 8.490 223.725 27.910 ;
        RECT 225.925 8.490 278.255 27.910 ;
        RECT 280.455 8.490 332.780 27.910 ;
        RECT 334.980 8.490 338.100 27.910 ;
  END
END N_term_single2
END LIBRARY

