VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO E_IO
  CLASS BLOCK ;
  FOREIGN E_IO ;
  ORIGIN 0.000 0.000 ;
  SIZE 110.000 BY 390.000 ;
  PIN A_I_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 1.400 110.000 1.960 ;
    END
  END A_I_top
  PIN A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 18.200 110.000 18.760 ;
    END
  END A_O_top
  PIN A_T_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 9.240 110.000 9.800 ;
    END
  END A_T_top
  PIN A_config_C_bit0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 51.800 110.000 52.360 ;
    END
  END A_config_C_bit0
  PIN A_config_C_bit1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 59.640 110.000 60.200 ;
    END
  END A_config_C_bit1
  PIN A_config_C_bit2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 68.600 110.000 69.160 ;
    END
  END A_config_C_bit2
  PIN A_config_C_bit3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 76.440 110.000 77.000 ;
    END
  END A_config_C_bit3
  PIN B_I_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 26.040 110.000 26.600 ;
    END
  END B_I_top
  PIN B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 42.840 110.000 43.400 ;
    END
  END B_O_top
  PIN B_T_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 35.000 110.000 35.560 ;
    END
  END B_T_top
  PIN B_config_C_bit0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 85.400 110.000 85.960 ;
    END
  END B_config_C_bit0
  PIN B_config_C_bit1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 93.240 110.000 93.800 ;
    END
  END B_config_C_bit1
  PIN B_config_C_bit2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 102.200 110.000 102.760 ;
    END
  END B_config_C_bit2
  PIN B_config_C_bit3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 111.160 110.000 111.720 ;
    END
  END B_config_C_bit3
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1.400 2.000 1.960 ;
    END
  END E1END[0]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3.640 2.000 4.200 ;
    END
  END E1END[1]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 7.000 2.000 7.560 ;
    END
  END E1END[2]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 10.360 2.000 10.920 ;
    END
  END E1END[3]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 37.240 2.000 37.800 ;
    END
  END E2END[0]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 40.600 2.000 41.160 ;
    END
  END E2END[1]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 42.840 2.000 43.400 ;
    END
  END E2END[2]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 46.200 2.000 46.760 ;
    END
  END E2END[3]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 49.560 2.000 50.120 ;
    END
  END E2END[4]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 52.920 2.000 53.480 ;
    END
  END E2END[5]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 55.160 2.000 55.720 ;
    END
  END E2END[6]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 58.520 2.000 59.080 ;
    END
  END E2END[7]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 12.600 2.000 13.160 ;
    END
  END E2MID[0]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 15.960 2.000 16.520 ;
    END
  END E2MID[1]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 19.320 2.000 19.880 ;
    END
  END E2MID[2]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 21.560 2.000 22.120 ;
    END
  END E2MID[3]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 24.920 2.000 25.480 ;
    END
  END E2MID[4]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 28.280 2.000 28.840 ;
    END
  END E2MID[5]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 31.640 2.000 32.200 ;
    END
  END E2MID[6]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 33.880 2.000 34.440 ;
    END
  END E2MID[7]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.040 2.000 110.600 ;
    END
  END E6END[0]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 140.280 2.000 140.840 ;
    END
  END E6END[10]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 143.640 2.000 144.200 ;
    END
  END E6END[11]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 113.400 2.000 113.960 ;
    END
  END E6END[1]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 116.760 2.000 117.320 ;
    END
  END E6END[2]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 119.000 2.000 119.560 ;
    END
  END E6END[3]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 122.360 2.000 122.920 ;
    END
  END E6END[4]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 125.720 2.000 126.280 ;
    END
  END E6END[5]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.960 2.000 128.520 ;
    END
  END E6END[6]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 131.320 2.000 131.880 ;
    END
  END E6END[7]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.680 2.000 135.240 ;
    END
  END E6END[8]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 136.920 2.000 137.480 ;
    END
  END E6END[9]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 61.880 2.000 62.440 ;
    END
  END EE4END[0]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 92.120 2.000 92.680 ;
    END
  END EE4END[10]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 95.480 2.000 96.040 ;
    END
  END EE4END[11]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 97.720 2.000 98.280 ;
    END
  END EE4END[12]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 101.080 2.000 101.640 ;
    END
  END EE4END[13]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 104.440 2.000 105.000 ;
    END
  END EE4END[14]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 106.680 2.000 107.240 ;
    END
  END EE4END[15]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 64.120 2.000 64.680 ;
    END
  END EE4END[1]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 67.480 2.000 68.040 ;
    END
  END EE4END[2]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.840 2.000 71.400 ;
    END
  END EE4END[3]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 74.200 2.000 74.760 ;
    END
  END EE4END[4]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 76.440 2.000 77.000 ;
    END
  END EE4END[5]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 79.800 2.000 80.360 ;
    END
  END EE4END[6]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 83.160 2.000 83.720 ;
    END
  END EE4END[7]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 85.400 2.000 85.960 ;
    END
  END EE4END[8]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 88.760 2.000 89.320 ;
    END
  END EE4END[9]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 292.600 2.000 293.160 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 322.840 2.000 323.400 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 326.200 2.000 326.760 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 328.440 2.000 329.000 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 331.800 2.000 332.360 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 335.160 2.000 335.720 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 337.400 2.000 337.960 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 340.760 2.000 341.320 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 344.120 2.000 344.680 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 347.480 2.000 348.040 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 349.720 2.000 350.280 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 294.840 2.000 295.400 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 353.080 2.000 353.640 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 356.440 2.000 357.000 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 358.680 2.000 359.240 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 362.040 2.000 362.600 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 365.400 2.000 365.960 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 368.760 2.000 369.320 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 371.000 2.000 371.560 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 374.360 2.000 374.920 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 377.720 2.000 378.280 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 379.960 2.000 380.520 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 298.200 2.000 298.760 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 383.320 2.000 383.880 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 386.680 2.000 387.240 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 301.560 2.000 302.120 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 304.920 2.000 305.480 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 307.160 2.000 307.720 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 310.520 2.000 311.080 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 313.880 2.000 314.440 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 316.120 2.000 316.680 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 319.480 2.000 320.040 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 119.000 110.000 119.560 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 204.120 110.000 204.680 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 211.960 110.000 212.520 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 220.920 110.000 221.480 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 228.760 110.000 229.320 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 237.720 110.000 238.280 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 245.560 110.000 246.120 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 254.520 110.000 255.080 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 262.360 110.000 262.920 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 271.320 110.000 271.880 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 279.160 110.000 279.720 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 127.960 110.000 128.520 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 288.120 110.000 288.680 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 297.080 110.000 297.640 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 304.920 110.000 305.480 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 313.880 110.000 314.440 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 321.720 110.000 322.280 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 330.680 110.000 331.240 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 338.520 110.000 339.080 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 347.480 110.000 348.040 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 355.320 110.000 355.880 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 364.280 110.000 364.840 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 135.800 110.000 136.360 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 372.120 110.000 372.680 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 381.080 110.000 381.640 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 144.760 110.000 145.320 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 152.600 110.000 153.160 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 161.560 110.000 162.120 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 169.400 110.000 169.960 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 178.360 110.000 178.920 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 186.200 110.000 186.760 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 195.160 110.000 195.720 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 5.880 0.000 6.440 2.000 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.400 0.000 57.960 2.000 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.000 0.000 63.560 2.000 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 68.600 0.000 69.160 2.000 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.080 0.000 73.640 2.000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 78.680 0.000 79.240 2.000 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 83.160 0.000 83.720 2.000 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 88.760 0.000 89.320 2.000 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.360 0.000 94.920 2.000 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 98.840 0.000 99.400 2.000 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.440 0.000 105.000 2.000 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 11.480 0.000 12.040 2.000 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 15.960 0.000 16.520 2.000 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 21.560 0.000 22.120 2.000 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 27.160 0.000 27.720 2.000 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 31.640 0.000 32.200 2.000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 37.240 0.000 37.800 2.000 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.720 0.000 42.280 2.000 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.320 0.000 47.880 2.000 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 52.920 0.000 53.480 2.000 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 5.880 388.000 6.440 390.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.400 388.000 57.960 390.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.000 388.000 63.560 390.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 68.600 388.000 69.160 390.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.080 388.000 73.640 390.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 78.680 388.000 79.240 390.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 83.160 388.000 83.720 390.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 88.760 388.000 89.320 390.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.360 388.000 94.920 390.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 98.840 388.000 99.400 390.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.440 388.000 105.000 390.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 11.480 388.000 12.040 390.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 15.960 388.000 16.520 390.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 21.560 388.000 22.120 390.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 27.160 388.000 27.720 390.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 31.640 388.000 32.200 390.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 37.240 388.000 37.800 390.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.720 388.000 42.280 390.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.320 388.000 47.880 390.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 52.920 388.000 53.480 390.000 ;
    END
  END FrameStrobe_O[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1.400 0.000 1.960 2.000 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1.400 388.000 1.960 390.000 ;
    END
  END UserCLKo
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 17.960 7.540 19.560 380.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 42.040 7.540 43.640 380.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 66.120 7.540 67.720 380.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 90.200 7.540 91.800 380.540 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 30.000 7.540 31.600 380.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 54.080 7.540 55.680 380.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 78.160 7.540 79.760 380.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 102.240 7.540 103.840 380.540 ;
    END
  END VSS
  PIN W1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 147.000 2.000 147.560 ;
    END
  END W1BEG[0]
  PIN W1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 149.240 2.000 149.800 ;
    END
  END W1BEG[1]
  PIN W1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 152.600 2.000 153.160 ;
    END
  END W1BEG[2]
  PIN W1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 155.960 2.000 156.520 ;
    END
  END W1BEG[3]
  PIN W2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 158.200 2.000 158.760 ;
    END
  END W2BEG[0]
  PIN W2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 161.560 2.000 162.120 ;
    END
  END W2BEG[1]
  PIN W2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.920 2.000 165.480 ;
    END
  END W2BEG[2]
  PIN W2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.280 2.000 168.840 ;
    END
  END W2BEG[3]
  PIN W2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 170.520 2.000 171.080 ;
    END
  END W2BEG[4]
  PIN W2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 173.880 2.000 174.440 ;
    END
  END W2BEG[5]
  PIN W2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 177.240 2.000 177.800 ;
    END
  END W2BEG[6]
  PIN W2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 179.480 2.000 180.040 ;
    END
  END W2BEG[7]
  PIN W2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.840 2.000 183.400 ;
    END
  END W2BEGb[0]
  PIN W2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 186.200 2.000 186.760 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 189.560 2.000 190.120 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 191.800 2.000 192.360 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 195.160 2.000 195.720 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.520 2.000 199.080 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 200.760 2.000 201.320 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 204.120 2.000 204.680 ;
    END
  END W2BEGb[7]
  PIN W6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 255.640 2.000 256.200 ;
    END
  END W6BEG[0]
  PIN W6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 285.880 2.000 286.440 ;
    END
  END W6BEG[10]
  PIN W6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 289.240 2.000 289.800 ;
    END
  END W6BEG[11]
  PIN W6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 259.000 2.000 259.560 ;
    END
  END W6BEG[1]
  PIN W6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.360 2.000 262.920 ;
    END
  END W6BEG[2]
  PIN W6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 264.600 2.000 265.160 ;
    END
  END W6BEG[3]
  PIN W6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 267.960 2.000 268.520 ;
    END
  END W6BEG[4]
  PIN W6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 271.320 2.000 271.880 ;
    END
  END W6BEG[5]
  PIN W6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 273.560 2.000 274.120 ;
    END
  END W6BEG[6]
  PIN W6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 276.920 2.000 277.480 ;
    END
  END W6BEG[7]
  PIN W6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 280.280 2.000 280.840 ;
    END
  END W6BEG[8]
  PIN W6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 283.640 2.000 284.200 ;
    END
  END W6BEG[9]
  PIN WW4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 207.480 2.000 208.040 ;
    END
  END WW4BEG[0]
  PIN WW4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 237.720 2.000 238.280 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 241.080 2.000 241.640 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 243.320 2.000 243.880 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 246.680 2.000 247.240 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 250.040 2.000 250.600 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 253.400 2.000 253.960 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 210.840 2.000 211.400 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 213.080 2.000 213.640 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 216.440 2.000 217.000 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 219.800 2.000 220.360 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 222.040 2.000 222.600 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 225.400 2.000 225.960 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 228.760 2.000 229.320 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 232.120 2.000 232.680 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 234.360 2.000 234.920 ;
    END
  END WW4BEG[9]
  OBS
      LAYER Metal1 ;
        RECT 6.720 7.540 103.840 380.540 ;
      LAYER Metal2 ;
        RECT 2.260 387.700 5.580 388.500 ;
        RECT 6.740 387.700 11.180 388.500 ;
        RECT 12.340 387.700 15.660 388.500 ;
        RECT 16.820 387.700 21.260 388.500 ;
        RECT 22.420 387.700 26.860 388.500 ;
        RECT 28.020 387.700 31.340 388.500 ;
        RECT 32.500 387.700 36.940 388.500 ;
        RECT 38.100 387.700 41.420 388.500 ;
        RECT 42.580 387.700 47.020 388.500 ;
        RECT 48.180 387.700 52.620 388.500 ;
        RECT 53.780 387.700 57.100 388.500 ;
        RECT 58.260 387.700 62.700 388.500 ;
        RECT 63.860 387.700 68.300 388.500 ;
        RECT 69.460 387.700 72.780 388.500 ;
        RECT 73.940 387.700 78.380 388.500 ;
        RECT 79.540 387.700 82.860 388.500 ;
        RECT 84.020 387.700 88.460 388.500 ;
        RECT 89.620 387.700 94.060 388.500 ;
        RECT 95.220 387.700 98.540 388.500 ;
        RECT 99.700 387.700 104.140 388.500 ;
        RECT 105.300 387.700 106.820 388.500 ;
        RECT 1.820 2.300 106.820 387.700 ;
        RECT 2.260 1.260 5.580 2.300 ;
        RECT 6.740 1.260 11.180 2.300 ;
        RECT 12.340 1.260 15.660 2.300 ;
        RECT 16.820 1.260 21.260 2.300 ;
        RECT 22.420 1.260 26.860 2.300 ;
        RECT 28.020 1.260 31.340 2.300 ;
        RECT 32.500 1.260 36.940 2.300 ;
        RECT 38.100 1.260 41.420 2.300 ;
        RECT 42.580 1.260 47.020 2.300 ;
        RECT 48.180 1.260 52.620 2.300 ;
        RECT 53.780 1.260 57.100 2.300 ;
        RECT 58.260 1.260 62.700 2.300 ;
        RECT 63.860 1.260 68.300 2.300 ;
        RECT 69.460 1.260 72.780 2.300 ;
        RECT 73.940 1.260 78.380 2.300 ;
        RECT 79.540 1.260 82.860 2.300 ;
        RECT 84.020 1.260 88.460 2.300 ;
        RECT 89.620 1.260 94.060 2.300 ;
        RECT 95.220 1.260 98.540 2.300 ;
        RECT 99.700 1.260 104.140 2.300 ;
        RECT 105.300 1.260 106.820 2.300 ;
      LAYER Metal3 ;
        RECT 2.300 386.380 108.500 386.820 ;
        RECT 1.260 384.180 108.500 386.380 ;
        RECT 2.300 383.020 108.500 384.180 ;
        RECT 1.260 381.940 108.500 383.020 ;
        RECT 1.260 380.820 107.700 381.940 ;
        RECT 2.300 380.780 107.700 380.820 ;
        RECT 2.300 379.660 108.500 380.780 ;
        RECT 1.260 378.580 108.500 379.660 ;
        RECT 2.300 377.420 108.500 378.580 ;
        RECT 1.260 375.220 108.500 377.420 ;
        RECT 2.300 374.060 108.500 375.220 ;
        RECT 1.260 372.980 108.500 374.060 ;
        RECT 1.260 371.860 107.700 372.980 ;
        RECT 2.300 371.820 107.700 371.860 ;
        RECT 2.300 370.700 108.500 371.820 ;
        RECT 1.260 369.620 108.500 370.700 ;
        RECT 2.300 368.460 108.500 369.620 ;
        RECT 1.260 366.260 108.500 368.460 ;
        RECT 2.300 365.140 108.500 366.260 ;
        RECT 2.300 365.100 107.700 365.140 ;
        RECT 1.260 363.980 107.700 365.100 ;
        RECT 1.260 362.900 108.500 363.980 ;
        RECT 2.300 361.740 108.500 362.900 ;
        RECT 1.260 359.540 108.500 361.740 ;
        RECT 2.300 358.380 108.500 359.540 ;
        RECT 1.260 357.300 108.500 358.380 ;
        RECT 2.300 356.180 108.500 357.300 ;
        RECT 2.300 356.140 107.700 356.180 ;
        RECT 1.260 355.020 107.700 356.140 ;
        RECT 1.260 353.940 108.500 355.020 ;
        RECT 2.300 352.780 108.500 353.940 ;
        RECT 1.260 350.580 108.500 352.780 ;
        RECT 2.300 349.420 108.500 350.580 ;
        RECT 1.260 348.340 108.500 349.420 ;
        RECT 2.300 347.180 107.700 348.340 ;
        RECT 1.260 344.980 108.500 347.180 ;
        RECT 2.300 343.820 108.500 344.980 ;
        RECT 1.260 341.620 108.500 343.820 ;
        RECT 2.300 340.460 108.500 341.620 ;
        RECT 1.260 339.380 108.500 340.460 ;
        RECT 1.260 338.260 107.700 339.380 ;
        RECT 2.300 338.220 107.700 338.260 ;
        RECT 2.300 337.100 108.500 338.220 ;
        RECT 1.260 336.020 108.500 337.100 ;
        RECT 2.300 334.860 108.500 336.020 ;
        RECT 1.260 332.660 108.500 334.860 ;
        RECT 2.300 331.540 108.500 332.660 ;
        RECT 2.300 331.500 107.700 331.540 ;
        RECT 1.260 330.380 107.700 331.500 ;
        RECT 1.260 329.300 108.500 330.380 ;
        RECT 2.300 328.140 108.500 329.300 ;
        RECT 1.260 327.060 108.500 328.140 ;
        RECT 2.300 325.900 108.500 327.060 ;
        RECT 1.260 323.700 108.500 325.900 ;
        RECT 2.300 322.580 108.500 323.700 ;
        RECT 2.300 322.540 107.700 322.580 ;
        RECT 1.260 321.420 107.700 322.540 ;
        RECT 1.260 320.340 108.500 321.420 ;
        RECT 2.300 319.180 108.500 320.340 ;
        RECT 1.260 316.980 108.500 319.180 ;
        RECT 2.300 315.820 108.500 316.980 ;
        RECT 1.260 314.740 108.500 315.820 ;
        RECT 2.300 313.580 107.700 314.740 ;
        RECT 1.260 311.380 108.500 313.580 ;
        RECT 2.300 310.220 108.500 311.380 ;
        RECT 1.260 308.020 108.500 310.220 ;
        RECT 2.300 306.860 108.500 308.020 ;
        RECT 1.260 305.780 108.500 306.860 ;
        RECT 2.300 304.620 107.700 305.780 ;
        RECT 1.260 302.420 108.500 304.620 ;
        RECT 2.300 301.260 108.500 302.420 ;
        RECT 1.260 299.060 108.500 301.260 ;
        RECT 2.300 297.940 108.500 299.060 ;
        RECT 2.300 297.900 107.700 297.940 ;
        RECT 1.260 296.780 107.700 297.900 ;
        RECT 1.260 295.700 108.500 296.780 ;
        RECT 2.300 294.540 108.500 295.700 ;
        RECT 1.260 293.460 108.500 294.540 ;
        RECT 2.300 292.300 108.500 293.460 ;
        RECT 1.260 290.100 108.500 292.300 ;
        RECT 2.300 288.980 108.500 290.100 ;
        RECT 2.300 288.940 107.700 288.980 ;
        RECT 1.260 287.820 107.700 288.940 ;
        RECT 1.260 286.740 108.500 287.820 ;
        RECT 2.300 285.580 108.500 286.740 ;
        RECT 1.260 284.500 108.500 285.580 ;
        RECT 2.300 283.340 108.500 284.500 ;
        RECT 1.260 281.140 108.500 283.340 ;
        RECT 2.300 280.020 108.500 281.140 ;
        RECT 2.300 279.980 107.700 280.020 ;
        RECT 1.260 278.860 107.700 279.980 ;
        RECT 1.260 277.780 108.500 278.860 ;
        RECT 2.300 276.620 108.500 277.780 ;
        RECT 1.260 274.420 108.500 276.620 ;
        RECT 2.300 273.260 108.500 274.420 ;
        RECT 1.260 272.180 108.500 273.260 ;
        RECT 2.300 271.020 107.700 272.180 ;
        RECT 1.260 268.820 108.500 271.020 ;
        RECT 2.300 267.660 108.500 268.820 ;
        RECT 1.260 265.460 108.500 267.660 ;
        RECT 2.300 264.300 108.500 265.460 ;
        RECT 1.260 263.220 108.500 264.300 ;
        RECT 2.300 262.060 107.700 263.220 ;
        RECT 1.260 259.860 108.500 262.060 ;
        RECT 2.300 258.700 108.500 259.860 ;
        RECT 1.260 256.500 108.500 258.700 ;
        RECT 2.300 255.380 108.500 256.500 ;
        RECT 2.300 255.340 107.700 255.380 ;
        RECT 1.260 254.260 107.700 255.340 ;
        RECT 2.300 254.220 107.700 254.260 ;
        RECT 2.300 253.100 108.500 254.220 ;
        RECT 1.260 250.900 108.500 253.100 ;
        RECT 2.300 249.740 108.500 250.900 ;
        RECT 1.260 247.540 108.500 249.740 ;
        RECT 2.300 246.420 108.500 247.540 ;
        RECT 2.300 246.380 107.700 246.420 ;
        RECT 1.260 245.260 107.700 246.380 ;
        RECT 1.260 244.180 108.500 245.260 ;
        RECT 2.300 243.020 108.500 244.180 ;
        RECT 1.260 241.940 108.500 243.020 ;
        RECT 2.300 240.780 108.500 241.940 ;
        RECT 1.260 238.580 108.500 240.780 ;
        RECT 2.300 237.420 107.700 238.580 ;
        RECT 1.260 235.220 108.500 237.420 ;
        RECT 2.300 234.060 108.500 235.220 ;
        RECT 1.260 232.980 108.500 234.060 ;
        RECT 2.300 231.820 108.500 232.980 ;
        RECT 1.260 229.620 108.500 231.820 ;
        RECT 2.300 228.460 107.700 229.620 ;
        RECT 1.260 226.260 108.500 228.460 ;
        RECT 2.300 225.100 108.500 226.260 ;
        RECT 1.260 222.900 108.500 225.100 ;
        RECT 2.300 221.780 108.500 222.900 ;
        RECT 2.300 221.740 107.700 221.780 ;
        RECT 1.260 220.660 107.700 221.740 ;
        RECT 2.300 220.620 107.700 220.660 ;
        RECT 2.300 219.500 108.500 220.620 ;
        RECT 1.260 217.300 108.500 219.500 ;
        RECT 2.300 216.140 108.500 217.300 ;
        RECT 1.260 213.940 108.500 216.140 ;
        RECT 2.300 212.820 108.500 213.940 ;
        RECT 2.300 212.780 107.700 212.820 ;
        RECT 1.260 211.700 107.700 212.780 ;
        RECT 2.300 211.660 107.700 211.700 ;
        RECT 2.300 210.540 108.500 211.660 ;
        RECT 1.260 208.340 108.500 210.540 ;
        RECT 2.300 207.180 108.500 208.340 ;
        RECT 1.260 204.980 108.500 207.180 ;
        RECT 2.300 203.820 107.700 204.980 ;
        RECT 1.260 201.620 108.500 203.820 ;
        RECT 2.300 200.460 108.500 201.620 ;
        RECT 1.260 199.380 108.500 200.460 ;
        RECT 2.300 198.220 108.500 199.380 ;
        RECT 1.260 196.020 108.500 198.220 ;
        RECT 2.300 194.860 107.700 196.020 ;
        RECT 1.260 192.660 108.500 194.860 ;
        RECT 2.300 191.500 108.500 192.660 ;
        RECT 1.260 190.420 108.500 191.500 ;
        RECT 2.300 189.260 108.500 190.420 ;
        RECT 1.260 187.060 108.500 189.260 ;
        RECT 2.300 185.900 107.700 187.060 ;
        RECT 1.260 183.700 108.500 185.900 ;
        RECT 2.300 182.540 108.500 183.700 ;
        RECT 1.260 180.340 108.500 182.540 ;
        RECT 2.300 179.220 108.500 180.340 ;
        RECT 2.300 179.180 107.700 179.220 ;
        RECT 1.260 178.100 107.700 179.180 ;
        RECT 2.300 178.060 107.700 178.100 ;
        RECT 2.300 176.940 108.500 178.060 ;
        RECT 1.260 174.740 108.500 176.940 ;
        RECT 2.300 173.580 108.500 174.740 ;
        RECT 1.260 171.380 108.500 173.580 ;
        RECT 2.300 170.260 108.500 171.380 ;
        RECT 2.300 170.220 107.700 170.260 ;
        RECT 1.260 169.140 107.700 170.220 ;
        RECT 2.300 169.100 107.700 169.140 ;
        RECT 2.300 167.980 108.500 169.100 ;
        RECT 1.260 165.780 108.500 167.980 ;
        RECT 2.300 164.620 108.500 165.780 ;
        RECT 1.260 162.420 108.500 164.620 ;
        RECT 2.300 161.260 107.700 162.420 ;
        RECT 1.260 159.060 108.500 161.260 ;
        RECT 2.300 157.900 108.500 159.060 ;
        RECT 1.260 156.820 108.500 157.900 ;
        RECT 2.300 155.660 108.500 156.820 ;
        RECT 1.260 153.460 108.500 155.660 ;
        RECT 2.300 152.300 107.700 153.460 ;
        RECT 1.260 150.100 108.500 152.300 ;
        RECT 2.300 148.940 108.500 150.100 ;
        RECT 1.260 147.860 108.500 148.940 ;
        RECT 2.300 146.700 108.500 147.860 ;
        RECT 1.260 145.620 108.500 146.700 ;
        RECT 1.260 144.500 107.700 145.620 ;
        RECT 2.300 144.460 107.700 144.500 ;
        RECT 2.300 143.340 108.500 144.460 ;
        RECT 1.260 141.140 108.500 143.340 ;
        RECT 2.300 139.980 108.500 141.140 ;
        RECT 1.260 137.780 108.500 139.980 ;
        RECT 2.300 136.660 108.500 137.780 ;
        RECT 2.300 136.620 107.700 136.660 ;
        RECT 1.260 135.540 107.700 136.620 ;
        RECT 2.300 135.500 107.700 135.540 ;
        RECT 2.300 134.380 108.500 135.500 ;
        RECT 1.260 132.180 108.500 134.380 ;
        RECT 2.300 131.020 108.500 132.180 ;
        RECT 1.260 128.820 108.500 131.020 ;
        RECT 2.300 127.660 107.700 128.820 ;
        RECT 1.260 126.580 108.500 127.660 ;
        RECT 2.300 125.420 108.500 126.580 ;
        RECT 1.260 123.220 108.500 125.420 ;
        RECT 2.300 122.060 108.500 123.220 ;
        RECT 1.260 119.860 108.500 122.060 ;
        RECT 2.300 118.700 107.700 119.860 ;
        RECT 1.260 117.620 108.500 118.700 ;
        RECT 2.300 116.460 108.500 117.620 ;
        RECT 1.260 114.260 108.500 116.460 ;
        RECT 2.300 113.100 108.500 114.260 ;
        RECT 1.260 112.020 108.500 113.100 ;
        RECT 1.260 110.900 107.700 112.020 ;
        RECT 2.300 110.860 107.700 110.900 ;
        RECT 2.300 109.740 108.500 110.860 ;
        RECT 1.260 107.540 108.500 109.740 ;
        RECT 2.300 106.380 108.500 107.540 ;
        RECT 1.260 105.300 108.500 106.380 ;
        RECT 2.300 104.140 108.500 105.300 ;
        RECT 1.260 103.060 108.500 104.140 ;
        RECT 1.260 101.940 107.700 103.060 ;
        RECT 2.300 101.900 107.700 101.940 ;
        RECT 2.300 100.780 108.500 101.900 ;
        RECT 1.260 98.580 108.500 100.780 ;
        RECT 2.300 97.420 108.500 98.580 ;
        RECT 1.260 96.340 108.500 97.420 ;
        RECT 2.300 95.180 108.500 96.340 ;
        RECT 1.260 94.100 108.500 95.180 ;
        RECT 1.260 92.980 107.700 94.100 ;
        RECT 2.300 92.940 107.700 92.980 ;
        RECT 2.300 91.820 108.500 92.940 ;
        RECT 1.260 89.620 108.500 91.820 ;
        RECT 2.300 88.460 108.500 89.620 ;
        RECT 1.260 86.260 108.500 88.460 ;
        RECT 2.300 85.100 107.700 86.260 ;
        RECT 1.260 84.020 108.500 85.100 ;
        RECT 2.300 82.860 108.500 84.020 ;
        RECT 1.260 80.660 108.500 82.860 ;
        RECT 2.300 79.500 108.500 80.660 ;
        RECT 1.260 77.300 108.500 79.500 ;
        RECT 2.300 76.140 107.700 77.300 ;
        RECT 1.260 75.060 108.500 76.140 ;
        RECT 2.300 73.900 108.500 75.060 ;
        RECT 1.260 71.700 108.500 73.900 ;
        RECT 2.300 70.540 108.500 71.700 ;
        RECT 1.260 69.460 108.500 70.540 ;
        RECT 1.260 68.340 107.700 69.460 ;
        RECT 2.300 68.300 107.700 68.340 ;
        RECT 2.300 67.180 108.500 68.300 ;
        RECT 1.260 64.980 108.500 67.180 ;
        RECT 2.300 63.820 108.500 64.980 ;
        RECT 1.260 62.740 108.500 63.820 ;
        RECT 2.300 61.580 108.500 62.740 ;
        RECT 1.260 60.500 108.500 61.580 ;
        RECT 1.260 59.380 107.700 60.500 ;
        RECT 2.300 59.340 107.700 59.380 ;
        RECT 2.300 58.220 108.500 59.340 ;
        RECT 1.260 56.020 108.500 58.220 ;
        RECT 2.300 54.860 108.500 56.020 ;
        RECT 1.260 53.780 108.500 54.860 ;
        RECT 2.300 52.660 108.500 53.780 ;
        RECT 2.300 52.620 107.700 52.660 ;
        RECT 1.260 51.500 107.700 52.620 ;
        RECT 1.260 50.420 108.500 51.500 ;
        RECT 2.300 49.260 108.500 50.420 ;
        RECT 1.260 47.060 108.500 49.260 ;
        RECT 2.300 45.900 108.500 47.060 ;
        RECT 1.260 43.700 108.500 45.900 ;
        RECT 2.300 42.540 107.700 43.700 ;
        RECT 1.260 41.460 108.500 42.540 ;
        RECT 2.300 40.300 108.500 41.460 ;
        RECT 1.260 38.100 108.500 40.300 ;
        RECT 2.300 36.940 108.500 38.100 ;
        RECT 1.260 35.860 108.500 36.940 ;
        RECT 1.260 34.740 107.700 35.860 ;
        RECT 2.300 34.700 107.700 34.740 ;
        RECT 2.300 33.580 108.500 34.700 ;
        RECT 1.260 32.500 108.500 33.580 ;
        RECT 2.300 31.340 108.500 32.500 ;
        RECT 1.260 29.140 108.500 31.340 ;
        RECT 2.300 27.980 108.500 29.140 ;
        RECT 1.260 26.900 108.500 27.980 ;
        RECT 1.260 25.780 107.700 26.900 ;
        RECT 2.300 25.740 107.700 25.780 ;
        RECT 2.300 24.620 108.500 25.740 ;
        RECT 1.260 22.420 108.500 24.620 ;
        RECT 2.300 21.260 108.500 22.420 ;
        RECT 1.260 20.180 108.500 21.260 ;
        RECT 2.300 19.060 108.500 20.180 ;
        RECT 2.300 19.020 107.700 19.060 ;
        RECT 1.260 17.900 107.700 19.020 ;
        RECT 1.260 16.820 108.500 17.900 ;
        RECT 2.300 15.660 108.500 16.820 ;
        RECT 1.260 13.460 108.500 15.660 ;
        RECT 2.300 12.300 108.500 13.460 ;
        RECT 1.260 11.220 108.500 12.300 ;
        RECT 2.300 10.100 108.500 11.220 ;
        RECT 2.300 10.060 107.700 10.100 ;
        RECT 1.260 8.940 107.700 10.060 ;
        RECT 1.260 7.860 108.500 8.940 ;
        RECT 2.300 6.700 108.500 7.860 ;
        RECT 1.260 4.500 108.500 6.700 ;
        RECT 2.300 3.340 108.500 4.500 ;
        RECT 1.260 2.260 108.500 3.340 ;
        RECT 2.300 1.820 107.700 2.260 ;
      LAYER Metal4 ;
        RECT 5.740 7.240 17.660 373.990 ;
        RECT 19.860 7.240 29.700 373.990 ;
        RECT 31.900 7.240 41.740 373.990 ;
        RECT 43.940 7.240 53.780 373.990 ;
        RECT 55.980 7.240 65.820 373.990 ;
        RECT 68.020 7.240 77.860 373.990 ;
        RECT 80.060 7.240 82.180 373.990 ;
        RECT 5.740 2.890 82.180 7.240 ;
  END
END E_IO
END LIBRARY

